module ORICDOS06
  (
   input wire [12:0] addr,
   input wire        clk,
   output logic [7:0]      data
   );

  logic [7:0]        rom_data[8192] =
    {8'h4c, 8'hc2, 8'he5, 8'h4c, 8'h0c, 8'he2, 8'h4c, 8'h34,
     8'heb, 8'h4c, 8'hce, 8'he4, 8'h4c, 8'hd3, 8'hea, 8'h4c,
     8'hde, 8'he4, 8'h4c, 8'hfc, 8'hea, 8'h4c, 8'h17, 8'he1,
     8'h4c, 8'h1f, 8'he1, 8'h4c, 8'hdc, 8'he7, 8'h4c, 8'h16,
     8'he8, 8'h4c, 8'h17, 8'he8, 8'h4c, 8'h25, 8'he8, 8'h4c,
     8'h2b, 8'he8, 8'h4c, 8'h46, 8'he8, 8'h4c, 8'h54, 8'he8,
     8'h4c, 8'h80, 8'he9, 8'h4c, 8'h72, 8'he8, 8'h4c, 8'h81,
     8'he8, 8'h4c, 8'h93, 8'he8, 8'h4c, 8'hb7, 8'he8, 8'h4c,
     8'hc5, 8'he8, 8'h4c, 8'hf6, 8'he8, 8'h4c, 8'h50, 8'he9,
     8'h4c, 8'ha8, 8'he9, 8'h4c, 8'hca, 8'he9, 8'h4c, 8'hb8,
     8'hea, 8'h4c, 8'hea, 8'hea, 8'h4c, 8'h27, 8'he1, 8'h4c,
     8'h2e, 8'he1, 8'h4c, 8'h70, 8'he0, 8'h4c, 8'h6a, 8'he1,
     8'h4c, 8'h63, 8'he1, 8'h4c, 8'hc7, 8'he4, 8'h4c, 8'h00,
     8'h00, 8'h4c, 8'h00, 8'h00, 8'h4c, 8'h45, 8'heb, 8'h00,
     8'h08, 8'h48, 8'h8a, 8'h48, 8'h98, 8'h48, 8'hba, 8'hbd,
     8'h05, 8'h01, 8'h18, 8'h85, 8'h0e, 8'h69, 8'h04, 8'h9d,
     8'h05, 8'h01, 8'hbd, 8'h06, 8'h01, 8'h85, 8'h0f, 8'h69,
     8'h00, 8'h9d, 8'h06, 8'h01, 8'ha0, 8'h01, 8'had, 8'h07,
     8'hc0, 8'hf0, 8'h02, 8'ha0, 8'h03, 8'hb1, 8'h0e, 8'h8d,
     8'h85, 8'h04, 8'hc8, 8'hb1, 8'h0e, 8'h8d, 8'h86, 8'h04,
     8'ha9, 8'h06, 8'h8d, 8'h81, 8'h04, 8'h68, 8'ha8, 8'h68,
     8'haa, 8'h68, 8'h28, 8'h4c, 8'h90, 8'h04, 8'h48, 8'had,
     8'h81, 8'h04, 8'h48, 8'had, 8'h85, 8'h04, 8'h48, 8'had,
     8'h86, 8'h04, 8'h48, 8'had, 8'h80, 8'h04, 8'h29, 8'hfe,
     8'h8d, 8'h80, 8'h04, 8'h8d, 8'h14, 8'h03, 8'ha9, 8'h00,
     8'h8d, 8'h85, 8'h04, 8'ha9, 8'h00, 8'h8d, 8'h86, 8'h04,
     8'ha9, 8'h06, 8'h8d, 8'h81, 8'h04, 8'h20, 8'h90, 8'h04,
     8'h68, 8'h8d, 8'h86, 8'h04, 8'h68, 8'h8d, 8'h85, 8'h04,
     8'h68, 8'h8d, 8'h81, 8'h04, 8'h68, 8'h40, 8'h48, 8'h8a,
     8'h48, 8'had, 8'h81, 8'h04, 8'h48, 8'had, 8'h85, 8'h04,
     8'h48, 8'had, 8'h86, 8'h04, 8'h48, 8'ha9, 8'h8a, 8'h8d,
     8'h85, 8'h04, 8'ha9, 8'h04, 8'h8d, 8'h86, 8'h04, 8'ha9,
     8'h06, 8'h8d, 8'h81, 8'h04, 8'h20, 8'h90, 8'h04, 8'h68,
     8'h8d, 8'h86, 8'h04, 8'h68, 8'h8d, 8'h85, 8'h04, 8'h68,
     8'h8d, 8'h81, 8'h04, 8'h68, 8'haa, 8'h68, 8'h40, 8'h20,
     8'h5a, 8'he0, 8'ha2, 8'hc5, 8'h92, 8'hc5, 8'h60, 8'h20,
     8'h5a, 8'he0, 8'hf8, 8'hc5, 8'he8, 8'hc5, 8'h60, 8'ha9,
     8'h0d, 8'h20, 8'h2e, 8'he1, 8'ha9, 8'h0a, 8'h08, 8'h8e,
     8'h51, 8'hc1, 8'haa, 8'h48, 8'ha5, 8'h0c, 8'h48, 8'ha5,
     8'h0d, 8'h48, 8'h20, 8'h5a, 8'he0, 8'h3f, 8'hf7, 8'h7c,
     8'hf7, 8'h68, 8'h85, 8'h0d, 8'h68, 8'h85, 8'h0c, 8'h68,
     8'hae, 8'h51, 8'hc1, 8'h28, 8'h60, 8'h48, 8'h4a, 8'h4a,
     8'h4a, 8'h4a, 8'h20, 8'h56, 8'he1, 8'h68, 8'h29, 8'h0f,
     8'h09, 8'h30, 8'hc9, 8'h3a, 8'h90, 8'hd0, 8'h69, 8'h06,
     8'hd0, 8'hcc, 8'hc8, 8'hb1, 8'he9, 8'hc9, 8'h20, 8'hf0,
     8'hf9, 8'h60, 8'ha9, 8'h00, 8'h8d, 8'h45, 8'hc1, 8'h8d,
     8'h46, 8'hc1, 8'hb1, 8'he9, 8'hc8, 8'hc9, 8'h20, 8'hf0,
     8'hf9, 8'hc9, 8'h23, 8'hd0, 8'h24, 8'hb1, 8'he9, 8'h20,
     8'hf1, 8'he1, 8'h90, 8'h1b, 8'hc8, 8'ha2, 8'h04, 8'h0e,
     8'h45, 8'hc1, 8'h2e, 8'h46, 8'hc1, 8'hca, 8'hd0, 8'hf7,
     8'h18, 8'h6d, 8'h45, 8'hc1, 8'h8d, 8'h45, 8'hc1, 8'h90,
     8'he4, 8'hee, 8'h46, 8'hc1, 8'h4c, 8'h7d, 8'he1, 8'h38,
     8'h60, 8'h88, 8'h20, 8'he6, 8'he1, 8'h90, 8'hf9, 8'hc8,
     8'h48, 8'had, 8'h46, 8'hc1, 8'h48, 8'had, 8'h45, 8'hc1,
     8'h0e, 8'h45, 8'hc1, 8'h2e, 8'h46, 8'hc1, 8'h0e, 8'h45,
     8'hc1, 8'h2e, 8'h46, 8'hc1, 8'h18, 8'h6d, 8'h45, 8'hc1,
     8'h8d, 8'h45, 8'hc1, 8'h68, 8'h6d, 8'h46, 8'hc1, 8'h8d,
     8'h46, 8'hc1, 8'h0e, 8'h45, 8'hc1, 8'h2e, 8'h46, 8'hc1,
     8'h68, 8'h18, 8'h6d, 8'h45, 8'hc1, 8'h8d, 8'h45, 8'hc1,
     8'h90, 8'h03, 8'hee, 8'h46, 8'hc1, 8'hb1, 8'he9, 8'h20,
     8'he6, 8'he1, 8'hb0, 8'hc3, 8'h38, 8'h60, 8'h38, 8'he9,
     8'h30, 8'h90, 8'h04, 8'hc9, 8'h0a, 8'h90, 8'hf5, 8'h18,
     8'h60, 8'h20, 8'he6, 8'he1, 8'hb0, 8'hee, 8'he9, 8'h06,
     8'hc9, 8'h10, 8'hb0, 8'hf3, 8'hc9, 8'h09, 8'h60, 8'h20,
     8'h5a, 8'he0, 8'ha3, 8'hc4, 8'h96, 8'hc4, 8'ha2, 8'ha0,
     8'hd0, 8'h02, 8'ha2, 8'h80, 8'h20, 8'he3, 8'he3, 8'h20,
     8'h1c, 8'he2, 8'h08, 8'h8a, 8'h48, 8'h20, 8'heb, 8'he3,
     8'h68, 8'haa, 8'h28, 8'h60, 8'h8e, 8'h05, 8'hc0, 8'h48,
     8'h98, 8'h48, 8'ha9, 8'h00, 8'h8d, 8'hfe, 8'h04, 8'ha9,
     8'h07, 8'h8d, 8'h08, 8'hc0, 8'h20, 8'ha2, 8'he2, 8'hf0,
     8'h16, 8'ha8, 8'h6a, 8'hb0, 8'h55, 8'ha9, 8'h20, 8'h2c,
     8'h05, 8'hc0, 8'h10, 8'h15, 8'h50, 8'h29, 8'hd0, 8'h4a,
     8'ha9, 8'h10, 8'h2c, 8'h05, 8'hc0, 8'hf0, 8'h3b, 8'ha2,
     8'h00, 8'h18, 8'h8e, 8'hfe, 8'h04, 8'h68, 8'ha8, 8'h68,
     8'h60, 8'h98, 8'h29, 8'h18, 8'hf0, 8'hf1, 8'hc0, 8'h18,
     8'hf0, 8'h30, 8'had, 8'h05, 8'hc0, 8'hc9, 8'h20, 8'hb0,
     8'h29, 8'hc9, 8'h10, 8'h90, 8'h1d, 8'hb0, 8'h10, 8'h98,
     8'h29, 8'h40, 8'hd0, 8'h1e, 8'hc0, 8'h10, 8'h90, 8'h12,
     8'had, 8'h05, 8'hc0, 8'h29, 8'h10, 8'hd0, 8'hd0, 8'hac,
     8'h05, 8'hc0, 8'h20, 8'h64, 8'he3, 8'h8c, 8'h05, 8'hc0,
     8'hb0, 8'h05, 8'hce, 8'h08, 8'hc0, 8'h10, 8'ha5, 8'h20,
     8'hb2, 8'he3, 8'ha2, 8'h01, 8'h38, 8'hb0, 8'hbe, 8'hc0,
     8'h20, 8'hb0, 8'h29, 8'hc0, 8'h10, 8'h90, 8'h25, 8'had,
     8'h01, 8'hc0, 8'h29, 8'h7f, 8'h8d, 8'h13, 8'h03, 8'h4c,
     8'hbc, 8'he2, 8'hac, 8'h05, 8'hc0, 8'h20, 8'h37, 8'he3,
     8'hb0, 8'h7b, 8'ha9, 8'h20, 8'h2c, 8'h05, 8'hc0, 8'h10,
     8'hde, 8'h50, 8'h10, 8'hd0, 8'h67, 8'ha9, 8'h10, 8'h2c,
     8'h05, 8'hc0, 8'hf0, 8'h2a, 8'h20, 8'h93, 8'he3, 8'h18,
     8'h58, 8'h90, 8'hfe, 8'had, 8'h01, 8'hc0, 8'h29, 8'h7f,
     8'hea, 8'hea, 8'hcd, 8'h11, 8'h03, 8'hf0, 8'h11, 8'had,
     8'h08, 8'hc0, 8'ha2, 8'h1c, 8'h20, 8'h1c, 8'he2, 8'h8d,
     8'h08, 8'hc0, 8'h8c, 8'h05, 8'hc0, 8'hb0, 8'h4e, 8'hea,
     8'had, 8'h02, 8'hc0, 8'h8d, 8'h12, 8'h03, 8'h98, 8'h29,
     8'h20, 8'hd0, 8'h1a, 8'h20, 8'h93, 8'he3, 8'h58, 8'had,
     8'h18, 8'h03, 8'h30, 8'hfb, 8'had, 8'h13, 8'h03, 8'h91,
     8'hfe, 8'hc8, 8'hd0, 8'hf3, 8'he6, 8'hff, 8'hd0, 8'hef,
     8'hf0, 8'h18, 8'hea, 8'hea, 8'hea, 8'h20, 8'h93, 8'he3,
     8'h58, 8'had, 8'h18, 8'h03, 8'h30, 8'hfb, 8'hb1, 8'hfe,
     8'h8d, 8'h13, 8'h03, 8'hc8, 8'hd0, 8'hf3, 8'he6, 8'hff,
     8'hd0, 8'hef, 8'hf0, 8'hfe, 8'had, 8'h05, 8'hc0, 8'h29,
     8'h10, 8'hf0, 8'hc8, 8'hd0, 8'he0, 8'h20, 8'hb2, 8'he3,
     8'had, 8'hfe, 8'h04, 8'h58, 8'h60, 8'had, 8'hfe, 8'h04,
     8'h29, 8'hbb, 8'h8d, 8'hfe, 8'h04, 8'h58, 8'h60, 8'had,
     8'h00, 8'hc0, 8'h29, 8'h03, 8'haa, 8'hbd, 8'hf3, 8'he3,
     8'h2c, 8'h01, 8'hc0, 8'h10, 8'h02, 8'h09, 8'h10, 8'h8d,
     8'h14, 8'h03, 8'haa, 8'had, 8'h80, 8'h04, 8'h8e, 8'h80,
     8'h04, 8'h29, 8'h7e, 8'h85, 8'hfe, 8'h8a, 8'h29, 8'h7e,
     8'hc5, 8'hfe, 8'hf0, 8'h31, 8'hc0, 8'h10, 8'h90, 8'h2d,
     8'hc0, 8'hf0, 8'hf0, 8'h29, 8'had, 8'h04, 8'hc0, 8'h48,
     8'ha9, 8'hc3, 8'h8d, 8'h04, 8'hc0, 8'had, 8'h08, 8'hc0,
     8'ha2, 8'hc0, 8'h20, 8'h1c, 8'he2, 8'h8d, 8'h08, 8'hc0,
     8'h68, 8'h8d, 8'h04, 8'hc0, 8'h8c, 8'h05, 8'hc0, 8'had,
     8'hfe, 8'h04, 8'hd0, 8'h0b, 8'had, 8'h12, 8'h03, 8'hea,
     8'hea, 8'hea, 8'h8d, 8'h11, 8'h03, 8'h18, 8'h60, 8'h38,
     8'h60, 8'hea, 8'hea, 8'h78, 8'h8c, 8'h05, 8'hc0, 8'had,
     8'h03, 8'hc0, 8'h85, 8'hfe, 8'had, 8'h04, 8'hc0, 8'h85,
     8'hff, 8'h8c, 8'h10, 8'h03, 8'had, 8'h80, 8'h04, 8'h09,
     8'h01, 8'h8d, 8'h14, 8'h03, 8'h8d, 8'h80, 8'h04, 8'ha0,
     8'h00, 8'h60, 8'had, 8'hfe, 8'h04, 8'ha2, 8'h08, 8'h20,
     8'h1c, 8'he2, 8'h8d, 8'hfe, 8'h04, 8'h60, 8'hea, 8'hea,
     8'h48, 8'had, 8'h14, 8'h03, 8'h30, 8'h19, 8'h68, 8'had,
     8'h80, 8'h04, 8'h29, 8'hfe, 8'h8d, 8'h80, 8'h04, 8'h8d,
     8'h14, 8'h03, 8'h68, 8'h68, 8'h68, 8'had, 8'h10, 8'h03,
     8'h29, 8'h5d, 8'h8d, 8'hfe, 8'h04, 8'h58, 8'h60, 8'h68,
     8'h4c, 8'he6, 8'he0, 8'h48, 8'ha9, 8'h40, 8'h8d, 8'h0e,
     8'h03, 8'h68, 8'h60, 8'h48, 8'ha9, 8'hc0, 8'h8d, 8'h0e,
     8'h03, 8'h68, 8'h60, 8'h04, 8'h24, 8'h44, 8'h64, 8'h20,
     8'h06, 8'he0, 8'h20, 8'h4b, 8'he0, 8'h20, 8'h45, 8'heb,
     8'h20, 8'h00, 8'he0, 8'h88, 8'hc8, 8'h20, 8'h60, 8'he0,
     8'h20, 8'h00, 8'h00, 8'hf0, 8'h55, 8'hc9, 8'h2c, 8'hd0,
     8'h15, 8'hc8, 8'hb1, 8'he9, 8'hc9, 8'h4e, 8'hd0, 8'h05,
     8'h8d, 8'h4f, 8'hc1, 8'h10, 8'he7, 8'hc9, 8'h44, 8'hd0,
     8'h0a, 8'h8d, 8'h50, 8'hc1, 8'h10, 8'hde, 8'ha2, 8'h01,
     8'h4c, 8'h1b, 8'he0, 8'hc9, 8'h4a, 8'hd0, 8'h15, 8'h8d,
     8'h41, 8'hc1, 8'ha5, 8'h9c, 8'h38, 8'he9, 8'h02, 8'h8d,
     8'h4d, 8'hc1, 8'ha5, 8'h9d, 8'he9, 8'h00, 8'h8d, 8'h4e,
     8'hc1, 8'h4c, 8'h04, 8'he4, 8'hc9, 8'h41, 8'hd0, 8'hde,
     8'h8d, 8'h4f, 8'hc1, 8'h8d, 8'h41, 8'hc1, 8'hc8, 8'h20,
     8'h5d, 8'he0, 8'h90, 8'hd2, 8'had, 8'h46, 8'hc1, 8'h8d,
     8'h4e, 8'hc1, 8'had, 8'h45, 8'hc1, 8'h8d, 8'h4d, 8'hc1,
     8'hb0, 8'ha3, 8'h98, 8'h48, 8'h20, 8'h09, 8'he0, 8'h68,
     8'ha8, 8'had, 8'h4c, 8'hc1, 8'hf0, 8'h08, 8'had, 8'h4f,
     8'hc1, 8'h10, 8'h03, 8'h6c, 8'h4b, 8'hc1, 8'had, 8'h4b,
     8'hc1, 8'hd0, 8'h03, 8'h4c, 8'h69, 8'he0, 8'hc9, 8'h03,
     8'hb0, 8'hf9, 8'h20, 8'h5a, 8'he0, 8'h6f, 8'hc5, 8'h5f,
     8'hc5, 8'ha5, 8'h92, 8'h85, 8'h9d, 8'h18, 8'ha5, 8'h91,
     8'h69, 8'h02, 8'h85, 8'h9c, 8'h90, 8'h02, 8'he6, 8'h9d,
     8'h85, 8'h9e, 8'h85, 8'ha0, 8'ha5, 8'h9d, 8'h85, 8'h9f,
     8'h85, 8'ha1, 8'ha5, 8'ha6, 8'h85, 8'ha2, 8'ha5, 8'ha7,
     8'h85, 8'ha3, 8'h20, 8'h5a, 8'he0, 8'h1f, 8'hc9, 8'h52,
     8'hc9, 8'h20, 8'h5a, 8'he0, 8'h65, 8'hc7, 8'h3a, 8'hc7,
     8'had, 8'h4b, 8'hc1, 8'hc9, 8'h01, 8'hf0, 8'h08, 8'h2c,
     8'h4f, 8'hc1, 8'h10, 8'h03, 8'h4c, 8'h69, 8'he0, 8'h20,
     8'h5a, 8'he0, 8'hb5, 8'hc4, 8'ha8, 8'hc4, 8'had, 8'h2b,
     8'hc1, 8'h8d, 8'h00, 8'hc0, 8'h20, 8'h2a, 8'he0, 8'h20,
     8'h0c, 8'he0, 8'he0, 8'h00, 8'hd0, 8'h05, 8'ha2, 8'h00,
     8'h4c, 8'h1b, 8'he0, 8'hbd, 8'h2f, 8'hc0, 8'h8d, 8'h01,
     8'hc0, 8'hbd, 8'h2e, 8'hc0, 8'h20, 8'h3f, 8'he8, 8'ha2,
     8'h00, 8'ha0, 8'h02, 8'h10, 8'h02, 8'h8a, 8'ha8, 8'had,
     8'h41, 8'hc1, 8'hd0, 8'h0c, 8'hb9, 8'h25, 8'hc0, 8'h8d,
     8'h4d, 8'hc1, 8'hb9, 8'h26, 8'hc0, 8'h8d, 8'h4e, 8'hc1,
     8'h38, 8'had, 8'h4d, 8'hc1, 8'hf9, 8'h25, 8'hc0, 8'h99,
     8'h25, 8'hc0, 8'had, 8'h4e, 8'hc1, 8'hf9, 8'h26, 8'hc0,
     8'h99, 8'h26, 8'hc0, 8'h18, 8'hb9, 8'h25, 8'hc0, 8'h79,
     8'h27, 8'hc0, 8'h99, 8'h27, 8'hc0, 8'hb9, 8'h26, 8'hc0,
     8'h79, 8'h28, 8'hc0, 8'h99, 8'h28, 8'hc0, 8'he0, 8'h00,
     8'hd0, 8'h0c, 8'hb9, 8'h2a, 8'hc0, 8'h8d, 8'h4c, 8'hc1,
     8'hb9, 8'h29, 8'hc0, 8'h8d, 8'h4b, 8'hc1, 8'had, 8'h50,
     8'hc1, 8'h30, 8'h36, 8'had, 8'h4e, 8'hc1, 8'h20, 8'h4d,
     8'he1, 8'had, 8'h4d, 8'hc1, 8'h20, 8'h4d, 8'he1, 8'ha9,
     8'h20, 8'h20, 8'h57, 8'he0, 8'hb9, 8'h28, 8'hc0, 8'h20,
     8'h4d, 8'he1, 8'hb9, 8'h27, 8'hc0, 8'h20, 8'h4d, 8'he1,
     8'had, 8'h41, 8'hc1, 8'hd0, 8'h11, 8'ha9, 8'h20, 8'h20,
     8'h57, 8'he0, 8'hb9, 8'h2a, 8'hc0, 8'h20, 8'h4d, 8'he1,
     8'hb9, 8'h29, 8'hc0, 8'h20, 8'h4d, 8'he1, 8'h20, 8'h54,
     8'he0, 8'had, 8'h4d, 8'hc1, 8'h85, 8'h0c, 8'had, 8'h4e,
     8'hc1, 8'h85, 8'h0d, 8'h18, 8'h98, 8'h69, 8'h08, 8'haa,
     8'hf0, 8'h25, 8'hbd, 8'h23, 8'hc0, 8'hf0, 8'h1d, 8'hc9,
     8'hff, 8'hd0, 8'h03, 8'h4c, 8'hf5, 8'he4, 8'h8d, 8'h41,
     8'hc1, 8'ha0, 8'h00, 8'he8, 8'hbd, 8'h23, 8'hc0, 8'h91,
     8'h0c, 8'he6, 8'h0c, 8'hd0, 8'h02, 8'he6, 8'h0d, 8'hce,
     8'h41, 8'hc1, 8'hd0, 8'hef, 8'he8, 8'hd0, 8'hdb, 8'had,
     8'h23, 8'hc0, 8'h8d, 8'h01, 8'hc0, 8'had, 8'h24, 8'hc0,
     8'hf0, 8'h07, 8'h20, 8'h3f, 8'he8, 8'ha2, 8'h02, 8'h10,
     8'hc9, 8'h60, 8'ha9, 8'hff, 8'h8d, 8'h4f, 8'hc1, 8'h8d,
     8'h50, 8'hc1, 8'h8d, 8'h3c, 8'hc1, 8'ha9, 8'h00, 8'h8d,
     8'h4d, 8'hc1, 8'h8d, 8'h4e, 8'hc1, 8'h8d, 8'h41, 8'hc1,
     8'h60, 8'h46, 8'h69, 8'h6c, 8'h65, 8'h20, 8'h6e, 8'h6f,
     8'h74, 8'h20, 8'h66, 8'h6f, 8'h75, 8'h6e, 8'h64, 8'h00,
     8'h49, 8'h6e, 8'h76, 8'h61, 8'h6c, 8'h69, 8'h64, 8'h20,
     8'h63, 8'h6f, 8'h6d, 8'h6d, 8'h61, 8'h6e, 8'h64, 8'h20,
     8'h65, 8'h6e, 8'h64, 8'h00, 8'h4e, 8'h6f, 8'h20, 8'h64,
     8'h72, 8'h69, 8'h76, 8'h65, 8'h20, 8'h6e, 8'h75, 8'h6d,
     8'h62, 8'h65, 8'h72, 8'h00, 8'h42, 8'h61, 8'h64, 8'h20,
     8'h64, 8'h72, 8'h69, 8'h76, 8'h65, 8'h20, 8'h6e, 8'h75,
     8'h6d, 8'h62, 8'h65, 8'h72, 8'h00, 8'h49, 8'h6e, 8'h76,
     8'h61, 8'h6c, 8'h69, 8'h64, 8'h20, 8'h66, 8'h69, 8'h6c,
     8'h65, 8'h6e, 8'h61, 8'h6d, 8'h65, 8'h00, 8'h44, 8'h69,
     8'h73, 8'h63, 8'h20, 8'h65, 8'h72, 8'h72, 8'h6f, 8'h72,
     8'h00, 8'h49, 8'h6c, 8'h6c, 8'h65, 8'h67, 8'h61, 8'h6c,
     8'h20, 8'h61, 8'h74, 8'h74, 8'h72, 8'h69, 8'h62, 8'h75,
     8'h74, 8'h65, 8'h00, 8'h57, 8'h69, 8'h6c, 8'h64, 8'h63,
     8'h61, 8'h72, 8'h64, 8'h28, 8'h73, 8'h29, 8'h20, 8'h6e,
     8'h6f, 8'h74, 8'h20, 8'h61, 8'h6c, 8'h6c, 8'h6f, 8'h77,
     8'h65, 8'h64, 8'h00, 8'h46, 8'h69, 8'h6c, 8'h65, 8'h20,
     8'h61, 8'h6c, 8'h72, 8'h65, 8'h61, 8'h64, 8'h79, 8'h20,
     8'h65, 8'h78, 8'h69, 8'h73, 8'h74, 8'h73, 8'h00, 8'h49,
     8'h6e, 8'h73, 8'h75, 8'h66, 8'h66, 8'h69, 8'h63, 8'h69,
     8'h65, 8'h6e, 8'h74, 8'h20, 8'h64, 8'h69, 8'h73, 8'h6b,
     8'h20, 8'h73, 8'h70, 8'h61, 8'h63, 8'h65, 8'h00, 8'h53,
     8'h74, 8'h61, 8'h72, 8'h74, 8'h20, 8'h61, 8'h64, 8'h64,
     8'h72, 8'h65, 8'h73, 8'h73, 8'h20, 8'h6d, 8'h69, 8'h73,
     8'h73, 8'h69, 8'h6e, 8'h67, 8'h00, 8'h49, 8'h6c, 8'h6c,
     8'h65, 8'h67, 8'h61, 8'h6c, 8'h20, 8'h71, 8'h75, 8'h61,
     8'h6e, 8'h74, 8'h69, 8'h74, 8'h79, 8'h00, 8'h45, 8'h6e,
     8'h64, 8'h20, 8'h61, 8'h64, 8'h64, 8'h72, 8'h65, 8'h73,
     8'h73, 8'h20, 8'h6d, 8'h69, 8'h73, 8'h73, 8'h69, 8'h6e,
     8'h67, 8'h00, 8'h53, 8'h74, 8'h61, 8'h72, 8'h74, 8'h20,
     8'h61, 8'h64, 8'h64, 8'h72, 8'h65, 8'h73, 8'h73, 8'h20,
     8'h3e, 8'h20, 8'h65, 8'h6e, 8'h64, 8'h20, 8'h61, 8'h64,
     8'h64, 8'h72, 8'h65, 8'h73, 8'h73, 8'h00, 8'h4d, 8'h69,
     8'h73, 8'h73, 8'h69, 8'h6e, 8'h67, 8'h20, 8'h27, 8'h54,
     8'h4f, 8'h27, 8'h00, 8'h52, 8'h65, 8'h6e, 8'h61, 8'h6d,
     8'h65, 8'h64, 8'h20, 8'h66, 8'h69, 8'h6c, 8'h65, 8'h20,
     8'h6e, 8'h6f, 8'h74, 8'h20, 8'h6f, 8'h6e, 8'h20, 8'h73,
     8'h61, 8'h6d, 8'h65, 8'h20, 8'h64, 8'h69, 8'h73, 8'h6b,
     8'h00, 8'h4d, 8'h69, 8'h73, 8'h73, 8'h69, 8'h6e, 8'h67,
     8'h20, 8'h63, 8'h6f, 8'h6d, 8'h6d, 8'h61, 8'h00, 8'h53,
     8'h6f, 8'h75, 8'h72, 8'h63, 8'h65, 8'h20, 8'h61, 8'h6e,
     8'h64, 8'h20, 8'h64, 8'h65, 8'h73, 8'h74, 8'h69, 8'h6e,
     8'h61, 8'h74, 8'h69, 8'h6f, 8'h6e, 8'h20, 8'h64, 8'h72,
     8'h69, 8'h76, 8'h65, 8'h73, 8'h20, 8'h6d, 8'h75, 8'h73,
     8'h74, 8'h20, 8'h62, 8'h65, 8'h20, 8'h73, 8'h61, 8'h6d,
     8'h65, 8'h00, 8'h44, 8'h65, 8'h73, 8'h74, 8'h69, 8'h6e,
     8'h61, 8'h74, 8'h69, 8'h6f, 8'h6e, 8'h20, 8'h6e, 8'h6f,
     8'h74, 8'h20, 8'h73, 8'h70, 8'h65, 8'h63, 8'h69, 8'h66,
     8'h69, 8'h65, 8'h64, 8'h00, 8'h43, 8'h61, 8'h6e, 8'h6e,
     8'h6f, 8'h74, 8'h20, 8'h6d, 8'h65, 8'h72, 8'h67, 8'h65,
     8'h20, 8'h61, 8'h6e, 8'h64, 8'h20, 8'h6f, 8'h76, 8'h65,
     8'h72, 8'h77, 8'h72, 8'h69, 8'h74, 8'h65, 8'h00, 8'h53,
     8'h69, 8'h6e, 8'h67, 8'h6c, 8'h65, 8'h20, 8'h64, 8'h65,
     8'h73, 8'h74, 8'h69, 8'h6e, 8'h61, 8'h74, 8'h69, 8'h6f,
     8'h6e, 8'h20, 8'h66, 8'h69, 8'h6c, 8'h65, 8'h20, 8'h6e,
     8'h6f, 8'h74, 8'h20, 8'h61, 8'h6c, 8'h6c, 8'h6f, 8'h77,
     8'h65, 8'h64, 8'h00, 8'h53, 8'h79, 8'h6e, 8'h74, 8'h61,
     8'h78, 8'h20, 8'h65, 8'h72, 8'h72, 8'h6f, 8'h72, 8'h00,
     8'hd9, 8'he8, 8'hfc, 8'h0c, 8'h1d, 8'h2e, 8'h39, 8'h4b,
     8'h63, 8'h77, 8'h8f, 8'ha5, 8'hb6, 8'hca, 8'he6, 8'hf3,
     8'h11, 8'h1f, 8'h4a, 8'h64, 8'h7f, 8'ha3, 8'he5, 8'he5,
     8'he5, 8'he6, 8'he6, 8'he6, 8'he6, 8'he6, 8'he6, 8'he6,
     8'he6, 8'he6, 8'he6, 8'he6, 8'he6, 8'he6, 8'he7, 8'he7,
     8'he7, 8'he7, 8'he7, 8'he7, 8'he8, 8'h8e, 8'hff, 8'h04,
     8'h6c, 8'h49, 8'hc1, 8'hca, 8'had, 8'hfd, 8'h04, 8'h29,
     8'h01, 8'hf0, 8'h03, 8'h4c, 8'h69, 8'he0, 8'he0, 8'h16,
     8'hb0, 8'h15, 8'hbd, 8'hb0, 8'he7, 8'h85, 8'h0c, 8'hbd,
     8'hc6, 8'he7, 8'h85, 8'h0d, 8'h20, 8'h2d, 8'he0, 8'ha9,
     8'h3a, 8'h20, 8'h57, 8'he0, 8'h4c, 8'h13, 8'he8, 8'h8a,
     8'h20, 8'h4d, 8'he1, 8'had, 8'hfe, 8'h04, 8'hf0, 8'h03,
     8'h20, 8'h4d, 8'he1, 8'h4c, 8'hff, 8'he1, 8'h60, 8'h20,
     8'h06, 8'he2, 8'had, 8'hfe, 8'h04, 8'hf0, 8'h05, 8'ha2,
     8'h05, 8'h4c, 8'h1b, 8'he0, 8'h60, 8'h20, 8'h0a, 8'he2,
     8'h4c, 8'h1a, 8'he8, 8'ha9, 8'h23, 8'h8d, 8'h03, 8'hc0,
     8'ha9, 8'hc0, 8'h8d, 8'h04, 8'hc0, 8'ha9, 8'h00, 8'h8d,
     8'h01, 8'hc0, 8'h8d, 8'h0a, 8'hc0, 8'ha9, 8'h01, 8'h8d,
     8'h02, 8'hc0, 8'h20, 8'h24, 8'he0, 8'h60, 8'hae, 8'h00,
     8'hc0, 8'hbd, 8'h13, 8'hc0, 8'hf0, 8'h01, 8'h60, 8'ha2,
     8'h03, 8'h4c, 8'h1b, 8'he0, 8'ha0, 8'h00, 8'hb1, 8'h0c,
     8'hf0, 8'h06, 8'h20, 8'h57, 8'he0, 8'hc8, 8'h10, 8'hf6,
     8'h60, 8'had, 8'h46, 8'hc1, 8'hd0, 8'h09, 8'had, 8'h45,
     8'hc1, 8'h30, 8'h04, 8'hc9, 8'h04, 8'h30, 8'h02, 8'ha9,
     8'hff, 8'h60, 8'h20, 8'h27, 8'he0, 8'ha2, 8'h07, 8'hbd,
     8'h33, 8'hc0, 8'h9d, 8'h23, 8'hc1, 8'hca, 8'h10, 8'hf7,
     8'h60, 8'h20, 8'h27, 8'he0, 8'ha2, 8'h07, 8'hbd, 8'h23,
     8'hc1, 8'h9d, 8'h33, 8'hc0, 8'hca, 8'h10, 8'hf7, 8'h20,
     8'h21, 8'he0, 8'h60, 8'had, 8'h3e, 8'hc1, 8'h8d, 8'h01,
     8'hc0, 8'had, 8'h3d, 8'hc1, 8'h20, 8'h3f, 8'he8, 8'ha2,
     8'h00, 8'hac, 8'h3f, 8'hc1, 8'hbd, 8'h2c, 8'hc1, 8'h99,
     8'h23, 8'hc0, 8'hc8, 8'he8, 8'he0, 8'h10, 8'hd0, 8'hf4,
     8'hee, 8'h25, 8'hc0, 8'h20, 8'h21, 8'he0, 8'h60, 8'h20,
     8'h3f, 8'he0, 8'hf0, 8'h08, 8'hee, 8'h29, 8'hc1, 8'hd0,
     8'h03, 8'hee, 8'h2a, 8'hc1, 8'h60, 8'had, 8'h23, 8'hc1,
     8'hf0, 8'h2b, 8'h8d, 8'h02, 8'hc0, 8'had, 8'h24, 8'hc1,
     8'h8d, 8'h01, 8'hc0, 8'h20, 8'h24, 8'he0, 8'had, 8'h24,
     8'hc0, 8'h8d, 8'h23, 8'hc1, 8'had, 8'h23, 8'hc0, 8'h8d,
     8'h24, 8'hc1, 8'h38, 8'had, 8'h27, 8'hc1, 8'he9, 8'h01,
     8'h8d, 8'h27, 8'hc1, 8'had, 8'h28, 8'hc1, 8'he9, 8'h00,
     8'h8d, 8'h28, 8'hc1, 8'ha9, 8'h01, 8'h60, 8'h20, 8'h24,
     8'he0, 8'had, 8'h25, 8'hc0, 8'hc9, 8'h0f, 8'hd0, 8'h31,
     8'had, 8'h24, 8'hc0, 8'hf0, 8'h0c, 8'h8d, 8'h02, 8'hc0,
     8'had, 8'h23, 8'hc0, 8'h8d, 8'h01, 8'hc0, 8'h4c, 8'hf6,
     8'he8, 8'had, 8'h23, 8'hc1, 8'hf0, 8'h39, 8'h8d, 8'h24,
     8'hc0, 8'had, 8'h24, 8'hc1, 8'h8d, 8'h23, 8'hc0, 8'h20,
     8'h21, 8'he0, 8'h20, 8'h3f, 8'he0, 8'ha9, 8'h00, 8'haa,
     8'h9d, 8'h23, 8'hc0, 8'he8, 8'hd0, 8'hfa, 8'h20, 8'h21,
     8'he0, 8'ha2, 8'h03, 8'hbd, 8'h23, 8'hc0, 8'hf0, 8'h07,
     8'h8a, 8'h18, 8'h69, 8'h10, 8'haa, 8'hd0, 8'hf4, 8'h8a,
     8'h8d, 8'h3f, 8'hc1, 8'had, 8'h01, 8'hc0, 8'h8d, 8'h3e,
     8'hc1, 8'had, 8'h02, 8'hc0, 8'h8d, 8'h3d, 8'hc1, 8'h60,
     8'h20, 8'h24, 8'he0, 8'hae, 8'h3f, 8'hc1, 8'hd0, 8'h28,
     8'h20, 8'h24, 8'he0, 8'ha2, 8'h03, 8'ha9, 8'h26, 8'h85,
     8'h0c, 8'ha9, 8'hc0, 8'h85, 8'h0d, 8'ha0, 8'h00, 8'hb1,
     8'h0c, 8'hf0, 8'h15, 8'ha0, 8'h08, 8'hb9, 8'h2c, 8'hc1,
     8'hc9, 8'h3f, 8'hf0, 8'h04, 8'hd1, 8'h0c, 8'hd0, 8'h08,
     8'h88, 8'h10, 8'hf2, 8'h8a, 8'h8d, 8'h3f, 8'hc1, 8'h60,
     8'h8a, 8'h18, 8'h69, 8'h10, 8'hb0, 8'h0e, 8'haa, 8'ha5,
     8'h0c, 8'h69, 8'h10, 8'h85, 8'h0c, 8'h90, 8'hd6, 8'he6,
     8'h0d, 8'h4c, 8'h65, 8'he9, 8'had, 8'h24, 8'hc0, 8'hf0,
     8'h0c, 8'h8d, 8'h02, 8'hc0, 8'had, 8'h23, 8'hc0, 8'h8d,
     8'h01, 8'hc0, 8'h4c, 8'h58, 8'he9, 8'ha2, 8'h00, 8'h60,
     8'had, 8'h13, 8'hc0, 8'hd0, 8'hfa, 8'h8d, 8'h00, 8'hc0,
     8'ha9, 8'h13, 8'h8d, 8'h03, 8'hc0, 8'ha9, 8'hc0, 8'h8d,
     8'h04, 8'hc0, 8'h4c, 8'h35, 8'he8, 8'h20, 8'h20, 8'h20,
     8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20, 8'h20,
     8'h20, 8'h00, 8'ha2, 8'h0b, 8'ha9, 8'h20, 8'h9d, 8'hbd,
     8'he9, 8'hca, 8'h10, 8'hfa, 8'h20, 8'h60, 8'he0, 8'h20,
     8'h00, 8'h00, 8'hf0, 8'h69, 8'h38, 8'he9, 8'h30, 8'hc9,
     8'h04, 8'hb0, 8'h0f, 8'hc8, 8'h8d, 8'h2b, 8'hc1, 8'ha2,
     8'h09, 8'ha9, 8'h20, 8'h9d, 8'h2b, 8'hc1, 8'hca, 8'hd0,
     8'hfa, 8'h60, 8'ha5, 8'hea, 8'h48, 8'ha5, 8'he9, 8'h48,
     8'h98, 8'h18, 8'h65, 8'he9, 8'h85, 8'he9, 8'h90, 8'h02,
     8'he6, 8'hea, 8'h20, 8'h5a, 8'he0, 8'h8b, 8'hce, 8'h17,
     8'hcf, 8'h24, 8'h28, 8'h10, 8'h56, 8'h20, 8'h5a, 8'he0,
     8'h15, 8'hd7, 8'hd0, 8'hd7, 8'hc9, 8'h0c, 8'h90, 8'h02,
     8'ha9, 8'h0c, 8'ha8, 8'h88, 8'h30, 8'h08, 8'hb1, 8'h91,
     8'h99, 8'hbd, 8'he9, 8'h4c, 8'h1b, 8'hea, 8'ha5, 8'he9,
     8'h48, 8'ha9, 8'hbd, 8'h85, 8'he9, 8'ha9, 8'he9, 8'h85,
     8'hea, 8'hc8, 8'h20, 8'h45, 8'hea, 8'h68, 8'h85, 8'hea,
     8'h68, 8'h18, 8'h85, 8'he9, 8'he5, 8'hea, 8'h49, 8'hff,
     8'ha8, 8'h68, 8'h85, 8'hea, 8'h60, 8'had, 8'h0c, 8'hc0,
     8'h8d, 8'h2b, 8'hc1, 8'h20, 8'he7, 8'he9, 8'hc8, 8'hb1,
     8'he9, 8'h88, 8'hc9, 8'hcd, 8'hf0, 8'h04, 8'hc9, 8'h2d,
     8'hd0, 8'h13, 8'hb1, 8'he9, 8'h38, 8'he9, 8'h30, 8'hc9,
     8'h04, 8'h90, 8'h05, 8'ha2, 8'h04, 8'h4c, 8'h1b, 8'he0,
     8'h8d, 8'h2b, 8'hc1, 8'hc8, 8'hc8, 8'ha2, 8'h00, 8'ha9,
     8'h06, 8'h20, 8'h8c, 8'hea, 8'hb1, 8'he9, 8'hc9, 8'h2e,
     8'hd0, 8'h08, 8'hc8, 8'ha2, 8'h06, 8'ha9, 8'h03, 8'h20,
     8'h8c, 8'hea, 8'h20, 8'h00, 8'h00, 8'hf0, 8'h04, 8'hc9,
     8'h20, 8'hd0, 8'hd8, 8'h60, 8'h8d, 8'h41, 8'hc1, 8'hb1,
     8'he9, 8'hc9, 8'h2a, 8'hf0, 8'h16, 8'hc9, 8'h3f, 8'hf0,
     8'h07, 8'h20, 8'h4e, 8'he0, 8'hc9, 8'h00, 8'hf0, 8'h0a,
     8'h9d, 8'h2c, 8'hc1, 8'he8, 8'hc8, 8'hce, 8'h41, 8'hc1,
     8'hd0, 8'he5, 8'h60, 8'ha9, 8'h3f, 8'h9d, 8'h2c, 8'hc1,
     8'he8, 8'hce, 8'h41, 8'hc1, 8'hd0, 8'hf7, 8'hc8, 8'h60,
     8'hc9, 8'h30, 8'h90, 8'h14, 8'hc9, 8'h3a, 8'h90, 8'h12,
     8'hc9, 8'h41, 8'h90, 8'h0c, 8'hc9, 8'h5b, 8'h90, 8'h0a,
     8'hc9, 8'h61, 8'h90, 8'h04, 8'hc9, 8'h7b, 8'h90, 8'h02,
     8'ha9, 8'h00, 8'h60, 8'h20, 8'h33, 8'he0, 8'had, 8'h26,
     8'hc1, 8'h8d, 8'h01, 8'hc0, 8'had, 8'h25, 8'hc1, 8'h8d,
     8'h02, 8'hc0, 8'ha9, 8'h00, 8'h8d, 8'h3f, 8'hc1, 8'h4c,
     8'h45, 8'he0, 8'ha2, 8'h09, 8'hac, 8'h3f, 8'hc1, 8'hb9,
     8'h2c, 8'hc0, 8'h9d, 8'h2c, 8'hc1, 8'hc8, 8'he8, 8'he0,
     8'h10, 8'hd0, 8'hf4, 8'h60, 8'hae, 8'h3f, 8'hc1, 8'ha0,
     8'h06, 8'hbd, 8'h23, 8'hc0, 8'hc9, 8'h20, 8'hd0, 8'h03,
     8'h20, 8'h57, 8'he0, 8'he8, 8'h88, 8'hd0, 8'hf2, 8'hae,
     8'h3f, 8'hc1, 8'ha0, 8'h06, 8'hbd, 8'h23, 8'hc0, 8'hc9,
     8'h20, 8'hf0, 8'h03, 8'h20, 8'h57, 8'he0, 8'he8, 8'h88,
     8'hd0, 8'hf2, 8'ha9, 8'h2e, 8'h20, 8'h57, 8'he0, 8'ha0,
     8'h03, 8'hbd, 8'h23, 8'hc0, 8'h20, 8'h57, 8'he0, 8'he8,
     8'h88, 8'hd0, 8'hf6, 8'h60, 8'ha5, 8'h0c, 8'h8d, 8'h47,
     8'hc1, 8'ha5, 8'h0d, 8'h8d, 8'h48, 8'hc1, 8'hba, 8'he8,
     8'he8, 8'h8e, 8'h40, 8'hc1, 8'h60, 8'ha2, 8'h08, 8'hbd,
     8'h2c, 8'hc1, 8'hc9, 8'h3f, 8'hf0, 8'h2b, 8'hca, 8'h10,
     8'hf6, 8'h60, 8'h43, 8'h4f, 8'h4d, 8'h20, 8'h06, 8'he0,
     8'ha0, 8'h00, 8'h98, 8'h20, 8'h48, 8'hea, 8'had, 8'h32,
     8'hc1, 8'hc9, 8'h20, 8'hd0, 8'h0b, 8'ha2, 8'h02, 8'hbd,
     8'h52, 8'heb, 8'h9d, 8'h32, 8'hc1, 8'hca, 8'h10, 8'hf7,
     8'h20, 8'h45, 8'heb, 8'h20, 8'h00, 8'he0, 8'h4c, 8'h62,
     8'he4, 8'ha2, 8'h07, 8'h4c, 8'h1b, 8'he0, 8'h78, 8'hd8,
     8'ha2, 8'hff, 8'h9a, 8'he8, 8'h8a, 8'ha8, 8'hca, 8'hd0,
     8'hfd, 8'h88, 8'hd0, 8'hfa, 8'h9d, 8'h00, 8'hc0, 8'h9d,
     8'h00, 8'hc1, 8'h95, 8'h00, 8'h9d, 8'h00, 8'h02, 8'hca,
     8'hd0, 8'hf2, 8'ha2, 8'h7a, 8'hbd, 8'hed, 8'hee, 8'h9d,
     8'h80, 8'h04, 8'hca, 8'h10, 8'hf7, 8'h20, 8'hae, 8'hee,
     8'ha2, 8'h0c, 8'hbd, 8'h68, 8'hef, 8'h9d, 8'he0, 8'hbf,
     8'hca, 8'h10, 8'hf7, 8'h20, 8'he0, 8'hbf, 8'hc0, 8'hea,
     8'hf0, 8'h0f, 8'ha9, 8'h01, 8'h8d, 8'h07, 8'hc0, 8'ha9,
     8'h44, 8'h8d, 8'hdc, 8'h04, 8'ha9, 8'h47, 8'h8d, 8'he4,
     8'h04, 8'ha2, 8'hff, 8'h86, 8'ha9, 8'ha9, 8'hff, 8'ha0,
     8'h97, 8'h85, 8'ha6, 8'h84, 8'ha7, 8'h8d, 8'hc1, 8'h02,
     8'h8c, 8'hc2, 8'h02, 8'h85, 8'ha2, 8'h84, 8'ha3, 8'ha2,
     8'h1c, 8'hbd, 8'hcf, 8'hee, 8'h95, 8'he1, 8'hca, 8'hd0,
     8'hf8, 8'had, 8'h07, 8'hc0, 8'hf0, 8'h28, 8'ha9, 8'hb9,
     8'h85, 8'hf0, 8'ha9, 8'hec, 8'h85, 8'hf1, 8'ha9, 8'h20,
     8'h8d, 8'h4e, 8'h02, 8'ha9, 8'h04, 8'h8d, 8'h4f, 8'h02,
     8'ha9, 8'h00, 8'h8d, 8'h60, 8'h02, 8'ha2, 8'h12, 8'hbd,
     8'h5d, 8'hee, 8'h9d, 8'h38, 8'h02, 8'hca, 8'h10, 8'hf7,
     8'ha9, 8'hb0, 8'ha0, 8'hcc, 8'h30, 8'h19, 8'ha9, 8'hff,
     8'ha0, 8'hbf, 8'h8d, 8'he1, 8'h02, 8'h8c, 8'he2, 8'h02,
     8'ha2, 8'h08, 8'hbd, 8'h54, 8'hee, 8'h9d, 8'h28, 8'h02,
     8'hca, 8'h10, 8'hf7, 8'ha9, 8'hed, 8'ha0, 8'hcb, 8'h85,
     8'h1b, 8'h84, 8'h1c, 8'ha9, 8'h4c, 8'h85, 8'h1a, 8'h85,
     8'hc3, 8'h85, 8'h21, 8'h8d, 8'hfb, 8'h02, 8'ha9, 8'ha0,
     8'ha0, 8'hd2, 8'hae, 8'h07, 8'hc0, 8'hf0, 8'h04, 8'ha9,
     8'h36, 8'ha0, 8'hd3, 8'h85, 8'h22, 8'h84, 8'h23, 8'h8d,
     8'hfc, 8'h02, 8'h8c, 8'hfd, 8'h02, 8'ha9, 8'hc4, 8'ha0,
     8'h04, 8'h8d, 8'hf5, 8'h02, 8'h8c, 8'hf6, 8'h02, 8'ha9,
     8'h00, 8'h8d, 8'hff, 8'h04, 8'h8d, 8'hfd, 8'h04, 8'h20,
     8'h5a, 8'he0, 8'h88, 8'hf8, 8'hb8, 8'hf8, 8'ha9, 8'h50,
     8'h85, 8'h31, 8'ha9, 8'h30, 8'h85, 8'h32, 8'ha9, 8'h03,
     8'h85, 8'hc2, 8'ha9, 8'h00, 8'h85, 8'hd7, 8'h85, 8'h88,
     8'h85, 8'h2f, 8'h48, 8'h8d, 8'h00, 8'h05, 8'h8d, 8'h01,
     8'h05, 8'h8d, 8'h02, 8'h05, 8'h8d, 8'hf7, 8'h02, 8'h85,
     8'h2e, 8'h8d, 8'hf1, 8'h02, 8'h8d, 8'hf2, 8'h02, 8'h8d,
     8'hf4, 8'h02, 8'ha9, 8'h88, 8'h85, 8'h85, 8'ha9, 8'h02,
     8'h8d, 8'hc0, 8'h02, 8'ha9, 8'h01, 8'ha0, 8'h05, 8'h85,
     8'h9a, 8'h84, 8'h9b, 8'ha9, 8'h03, 8'h85, 8'h9c, 8'h84,
     8'h9d, 8'h85, 8'h9e, 8'h84, 8'h9f, 8'h85, 8'ha0, 8'h84,
     8'ha1, 8'ha2, 8'h00, 8'h20, 8'h92, 8'hee, 8'ha2, 8'h09,
     8'hbd, 8'h40, 8'hee, 8'h9d, 8'h2b, 8'hc1, 8'hca, 8'h10,
     8'hf7, 8'ha9, 8'h8a, 8'h8d, 8'h49, 8'hc1, 8'ha9, 8'hee,
     8'h8d, 8'h4a, 8'hc1, 8'ha2, 8'hd8, 8'h8e, 8'h10, 8'h03,
     8'ha2, 8'h08, 8'h20, 8'h03, 8'he0, 8'h20, 8'h48, 8'he0,
     8'h20, 8'h00, 8'he0, 8'h20, 8'h09, 8'he0, 8'h20, 8'ha3,
     8'hee, 8'ha2, 8'h08, 8'hbd, 8'h5a, 8'hed, 8'h95, 8'h35,
     8'hca, 8'h10, 8'hf8, 8'ha2, 8'hff, 8'he8, 8'hbd, 8'hd0,
     8'h9f, 8'h9d, 8'h82, 8'hbb, 8'hd0, 8'hf7, 8'ha2, 8'h1a,
     8'hbd, 8'h3f, 8'hed, 8'h9d, 8'he0, 8'hbf, 8'hca, 8'h10,
     8'hf7, 8'ha9, 8'hae, 8'ha0, 8'hed, 8'hae, 8'h07, 8'hc0,
     8'hf0, 8'h04, 8'ha9, 8'hf1, 8'ha0, 8'hed, 8'h85, 8'h0c,
     8'h84, 8'h0d, 8'h20, 8'h2d, 8'he0, 8'ha2, 8'h09, 8'hbd,
     8'h4a, 8'hee, 8'h9d, 8'h2b, 8'hc1, 8'hca, 8'h10, 8'hf7,
     8'h20, 8'h0c, 8'he0, 8'he0, 8'h00, 8'hd0, 8'h0d, 8'h86,
     8'h35, 8'ha9, 8'h35, 8'h85, 8'h0c, 8'ha9, 8'hee, 8'h85,
     8'h0d, 8'h20, 8'h2d, 8'he0, 8'h4c, 8'he0, 8'hbf, 8'h78,
     8'ha9, 8'h84, 8'h8d, 8'h80, 8'h04, 8'h8d, 8'h14, 8'h03,
     8'h20, 8'hf8, 8'hbf, 8'ha2, 8'h34, 8'ha0, 8'h00, 8'h58,
     8'h20, 8'h5a, 8'hd4, 8'hcd, 8'hc4, 8'hbd, 8'hc4, 8'h6c,
     8'h4b, 8'hc1, 8'h21, 8'h42, 8'h4f, 8'h4f, 8'h54, 8'h55,
     8'h50, 8'h00, 8'h00, 8'h69, 8'h6e, 8'h73, 8'h65, 8'h72,
     8'h74, 8'h20, 8'h73, 8'h79, 8'h73, 8'h74, 8'h65, 8'h6d,
     8'h20, 8'h64, 8'h69, 8'h73, 8'h63, 8'h00, 8'h0c, 8'h4e,
     8'h6f, 8'h20, 8'h6f, 8'h70, 8'h65, 8'h72, 8'h61, 8'h74,
     8'h69, 8'h6e, 8'h67, 8'h20, 8'h73, 8'h79, 8'h73, 8'h74,
     8'h65, 8'h6d, 8'h20, 8'h6f, 8'h6e, 8'h20, 8'h64, 8'h69,
     8'h73, 8'h63, 8'h08, 8'h00, 8'h0c, 8'h52, 8'h56, 8'h31,
     8'h20, 8'h61, 8'h64, 8'h6a, 8'h75, 8'h73, 8'h74, 8'h6d,
     8'h65, 8'h6e, 8'h74, 8'h20, 8'h72, 8'h65, 8'h71, 8'h75,
     8'h69, 8'h72, 8'h65, 8'h64, 8'h08, 8'h00, 8'h0c, 8'h4f,
     8'h52, 8'h49, 8'h43, 8'h20, 8'h45, 8'h58, 8'h54, 8'h45,
     8'h4e, 8'h44, 8'h45, 8'h44, 8'h20, 8'h42, 8'h41, 8'h53,
     8'h49, 8'h43, 8'h20, 8'h56, 8'h31, 8'h2e, 8'h30, 8'h0d,
     8'h0a, 8'h60, 8'h20, 8'h31, 8'h39, 8'h38, 8'h33, 8'h20,
     8'h54, 8'h41, 8'h4e, 8'h47, 8'h45, 8'h52, 8'h49, 8'h4e,
     8'h45, 8'h0d, 8'h0a, 8'h0a, 8'h0a, 8'h34, 8'h37, 8'h38,
     8'h37, 8'h30, 8'h20, 8'h42, 8'h59, 8'h54, 8'h45, 8'h53,
     8'h20, 8'h46, 8'h52, 8'h45, 8'h45, 8'h0d, 8'h0a, 8'h0a,
     8'h00, 8'h0c, 8'h4f, 8'h52, 8'h49, 8'h43, 8'h20, 8'h45,
     8'h58, 8'h54, 8'h45, 8'h4e, 8'h44, 8'h45, 8'h44, 8'h20,
     8'h42, 8'h41, 8'h53, 8'h49, 8'h43, 8'h20, 8'h56, 8'h31,
     8'h2e, 8'h31, 8'h0d, 8'h0a, 8'h60, 8'h20, 8'h31, 8'h39,
     8'h38, 8'h33, 8'h20, 8'h54, 8'h41, 8'h4e, 8'h47, 8'h45,
     8'h52, 8'h49, 8'h4e, 8'h45, 8'h0d, 8'h0a, 8'h0a, 8'h0a,
     8'h20, 8'h33, 8'h37, 8'h36, 8'h33, 8'h31, 8'h20, 8'h42,
     8'h59, 8'h54, 8'h45, 8'h53, 8'h20, 8'h46, 8'h52, 8'h45,
     8'h45, 8'h0d, 8'h0a, 8'h0a, 8'h00, 8'h0d, 8'h0a, 8'h52,
     8'h65, 8'h61, 8'h64, 8'h79, 8'h20, 8'h0d, 8'h0a, 8'h00,
     8'h00, 8'h53, 8'h59, 8'h53, 8'h54, 8'h45, 8'h4d, 8'h44,
     8'h4f, 8'h53, 8'h00, 8'h42, 8'h4f, 8'h4f, 8'h54, 8'h55,
     8'h50, 8'h43, 8'h4f, 8'h4d, 8'h4c, 8'h03, 8'hec, 8'h4c,
     8'h30, 8'hf4, 8'h01, 8'h00, 8'h40, 8'h4c, 8'h7c, 8'hf7,
     8'h4c, 8'h78, 8'heb, 8'h4c, 8'hc1, 8'hf5, 8'h4c, 8'h65,
     8'hf8, 8'h4c, 8'h22, 8'hee, 8'h4c, 8'hb2, 8'hf8, 8'h40,
     8'ha2, 8'h31, 8'ha0, 8'h00, 8'ha9, 8'h1a, 8'h99, 8'h80,
     8'hbb, 8'h99, 8'h80, 8'hbc, 8'h99, 8'h80, 8'hbd, 8'h99,
     8'h80, 8'hbe, 8'h99, 8'hfe, 8'hbe, 8'h88, 8'hd0, 8'hee,
     8'hf0, 8'h02, 8'ha2, 8'h13, 8'h20, 8'h92, 8'hee, 8'h4c,
     8'h8f, 8'hee, 8'h20, 8'ha3, 8'hee, 8'h4c, 8'h9d, 8'hee,
     8'he8, 8'h99, 8'h82, 8'hbb, 8'hc8, 8'hbd, 8'h63, 8'hed,
     8'hd0, 8'hf6, 8'h60, 8'ha0, 8'h1b, 8'ha9, 8'h20, 8'h99,
     8'h81, 8'hbb, 8'h88, 8'hd0, 8'hfa, 8'h60, 8'ha2, 8'h00,
     8'hbd, 8'ha5, 8'hc0, 8'ha8, 8'ha9, 8'h55, 8'h9d, 8'ha5,
     8'hc0, 8'hdd, 8'ha5, 8'hc0, 8'hd0, 8'hb2, 8'ha9, 8'haa,
     8'h9d, 8'ha5, 8'hc0, 8'hdd, 8'ha5, 8'hc0, 8'hd0, 8'ha8,
     8'h98, 8'h9d, 8'ha5, 8'hc0, 8'he8, 8'hd0, 8'he1, 8'h60,
     8'he6, 8'he9, 8'hd0, 8'h02, 8'he6, 8'hea, 8'had, 8'h60,
     8'hea, 8'hc9, 8'h20, 8'hf0, 8'hf3, 8'h20, 8'h41, 8'hea,
     8'h60, 8'h2c, 8'h60, 8'hea, 8'h2c, 8'h60, 8'hea, 8'h60,
     8'h80, 8'h4f, 8'hc7, 8'h52, 8'h58, 8'h04, 8'h00, 8'h00,
     8'h00, 8'h4c, 8'h60, 8'hea, 8'h4c, 8'he6, 8'h04, 8'h4c,
     8'hd6, 8'h04, 8'h4c, 8'hde, 8'h04, 8'h08, 8'h78, 8'h8d,
     8'h82, 8'h04, 8'h68, 8'h8d, 8'h83, 8'h04, 8'had, 8'h80,
     8'h04, 8'h48, 8'had, 8'h81, 8'h04, 8'h20, 8'he6, 8'h04,
     8'had, 8'h83, 8'h04, 8'h48, 8'had, 8'h82, 8'h04, 8'h28,
     8'h20, 8'h84, 8'h04, 8'h08, 8'h78, 8'h8d, 8'h82, 8'h04,
     8'h68, 8'h8d, 8'h83, 8'h04, 8'h68, 8'h20, 8'he6, 8'h04,
     8'had, 8'h83, 8'h04, 8'h48, 8'had, 8'h82, 8'h04, 8'h28,
     8'h60, 8'ha9, 8'h00, 8'h8d, 8'h81, 8'h04, 8'ha9, 8'h66,
     8'h8d, 8'h85, 8'h04, 8'ha9, 8'hd4, 8'h8d, 8'h86, 8'h04,
     8'h4c, 8'h90, 8'h04, 8'h08, 8'hba, 8'hfe, 8'h02, 8'h01,
     8'h4c, 8'h28, 8'h02, 8'h08, 8'hba, 8'hfe, 8'h02, 8'h01,
     8'h4c, 8'h2b, 8'h02, 8'h78, 8'h29, 8'h02, 8'h8d, 8'h81,
     8'h04, 8'had, 8'h80, 8'h04, 8'h29, 8'hfd, 8'h0d, 8'h81,
     8'h04, 8'h8d, 8'h14, 8'h03, 8'h8d, 8'h80, 8'h04, 8'h60,
     8'ha9, 8'h06, 8'h20, 8'h87, 8'h04, 8'hac, 8'h02, 8'hc0,
     8'ha9, 8'h00, 8'h4c, 8'h87, 8'h04, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff, 8'hff,
     8'h4f, 8'h72, 8'h69, 8'h63, 8'h20, 8'h44, 8'h4f, 8'h53,
     8'h20, 8'h56, 8'h30, 8'h2e, 8'h36, 8'h00, 8'h00, 8'h00,
     8'h28, 8'h43, 8'h29, 8'h20, 8'h4f, 8'h52, 8'h49, 8'h43,
     8'h20, 8'h31, 8'h39, 8'h38, 8'h33, 8'h00, 8'h00, 8'h00,
     8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00, 8'h00,
     8'h00, 8'h00, 8'hae, 8'he0, 8'h7e, 8'heb, 8'hc0, 8'he3};

  always @(posedge clk) begin
    data <= rom_data[addr];
  end
endmodule // ORICDOS06
