library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ORICDOS06VHDL is
 port (
   addr : in  std_logic_vector( 12 downto 0);
   clk  : in  std_logic;
   data : out std_logic_vector(7 downto 0)
   );
end entity;

architecture prom of ORICDOS06VHDL is
  type rom is array(0 to 8191) of std_logic_vector(7 downto 0);
  signal rom_data: rom := (
     X"4c", X"c2", X"e5", X"4c", X"0c", X"e2", X"4c", X"34",
     X"eb", X"4c", X"ce", X"e4", X"4c", X"d3", X"ea", X"4c",
     X"de", X"e4", X"4c", X"fc", X"ea", X"4c", X"17", X"e1",
     X"4c", X"1f", X"e1", X"4c", X"dc", X"e7", X"4c", X"16",
     X"e8", X"4c", X"17", X"e8", X"4c", X"25", X"e8", X"4c",
     X"2b", X"e8", X"4c", X"46", X"e8", X"4c", X"54", X"e8",
     X"4c", X"80", X"e9", X"4c", X"72", X"e8", X"4c", X"81",
     X"e8", X"4c", X"93", X"e8", X"4c", X"b7", X"e8", X"4c",
     X"c5", X"e8", X"4c", X"f6", X"e8", X"4c", X"50", X"e9",
     X"4c", X"a8", X"e9", X"4c", X"ca", X"e9", X"4c", X"b8",
     X"ea", X"4c", X"ea", X"ea", X"4c", X"27", X"e1", X"4c",
     X"2e", X"e1", X"4c", X"70", X"e0", X"4c", X"6a", X"e1",
     X"4c", X"63", X"e1", X"4c", X"c7", X"e4", X"4c", X"00",
     X"00", X"4c", X"00", X"00", X"4c", X"45", X"eb", X"00",
     X"08", X"48", X"8a", X"48", X"98", X"48", X"ba", X"bd",
     X"05", X"01", X"18", X"85", X"0e", X"69", X"04", X"9d",
     X"05", X"01", X"bd", X"06", X"01", X"85", X"0f", X"69",
     X"00", X"9d", X"06", X"01", X"a0", X"01", X"ad", X"07",
     X"c0", X"f0", X"02", X"a0", X"03", X"b1", X"0e", X"8d",
     X"85", X"04", X"c8", X"b1", X"0e", X"8d", X"86", X"04",
     X"a9", X"06", X"8d", X"81", X"04", X"68", X"a8", X"68",
     X"aa", X"68", X"28", X"4c", X"90", X"04", X"48", X"ad",
     X"81", X"04", X"48", X"ad", X"85", X"04", X"48", X"ad",
     X"86", X"04", X"48", X"ad", X"80", X"04", X"29", X"fe",
     X"8d", X"80", X"04", X"8d", X"14", X"03", X"a9", X"00",
     X"8d", X"85", X"04", X"a9", X"00", X"8d", X"86", X"04",
     X"a9", X"06", X"8d", X"81", X"04", X"20", X"90", X"04",
     X"68", X"8d", X"86", X"04", X"68", X"8d", X"85", X"04",
     X"68", X"8d", X"81", X"04", X"68", X"40", X"48", X"8a",
     X"48", X"ad", X"81", X"04", X"48", X"ad", X"85", X"04",
     X"48", X"ad", X"86", X"04", X"48", X"a9", X"8a", X"8d",
     X"85", X"04", X"a9", X"04", X"8d", X"86", X"04", X"a9",
     X"06", X"8d", X"81", X"04", X"20", X"90", X"04", X"68",
     X"8d", X"86", X"04", X"68", X"8d", X"85", X"04", X"68",
     X"8d", X"81", X"04", X"68", X"aa", X"68", X"40", X"20",
     X"5a", X"e0", X"a2", X"c5", X"92", X"c5", X"60", X"20",
     X"5a", X"e0", X"f8", X"c5", X"e8", X"c5", X"60", X"a9",
     X"0d", X"20", X"2e", X"e1", X"a9", X"0a", X"08", X"8e",
     X"51", X"c1", X"aa", X"48", X"a5", X"0c", X"48", X"a5",
     X"0d", X"48", X"20", X"5a", X"e0", X"3f", X"f7", X"7c",
     X"f7", X"68", X"85", X"0d", X"68", X"85", X"0c", X"68",
     X"ae", X"51", X"c1", X"28", X"60", X"48", X"4a", X"4a",
     X"4a", X"4a", X"20", X"56", X"e1", X"68", X"29", X"0f",
     X"09", X"30", X"c9", X"3a", X"90", X"d0", X"69", X"06",
     X"d0", X"cc", X"c8", X"b1", X"e9", X"c9", X"20", X"f0",
     X"f9", X"60", X"a9", X"00", X"8d", X"45", X"c1", X"8d",
     X"46", X"c1", X"b1", X"e9", X"c8", X"c9", X"20", X"f0",
     X"f9", X"c9", X"23", X"d0", X"24", X"b1", X"e9", X"20",
     X"f1", X"e1", X"90", X"1b", X"c8", X"a2", X"04", X"0e",
     X"45", X"c1", X"2e", X"46", X"c1", X"ca", X"d0", X"f7",
     X"18", X"6d", X"45", X"c1", X"8d", X"45", X"c1", X"90",
     X"e4", X"ee", X"46", X"c1", X"4c", X"7d", X"e1", X"38",
     X"60", X"88", X"20", X"e6", X"e1", X"90", X"f9", X"c8",
     X"48", X"ad", X"46", X"c1", X"48", X"ad", X"45", X"c1",
     X"0e", X"45", X"c1", X"2e", X"46", X"c1", X"0e", X"45",
     X"c1", X"2e", X"46", X"c1", X"18", X"6d", X"45", X"c1",
     X"8d", X"45", X"c1", X"68", X"6d", X"46", X"c1", X"8d",
     X"46", X"c1", X"0e", X"45", X"c1", X"2e", X"46", X"c1",
     X"68", X"18", X"6d", X"45", X"c1", X"8d", X"45", X"c1",
     X"90", X"03", X"ee", X"46", X"c1", X"b1", X"e9", X"20",
     X"e6", X"e1", X"b0", X"c3", X"38", X"60", X"38", X"e9",
     X"30", X"90", X"04", X"c9", X"0a", X"90", X"f5", X"18",
     X"60", X"20", X"e6", X"e1", X"b0", X"ee", X"e9", X"06",
     X"c9", X"10", X"b0", X"f3", X"c9", X"09", X"60", X"20",
     X"5a", X"e0", X"a3", X"c4", X"96", X"c4", X"a2", X"a0",
     X"d0", X"02", X"a2", X"80", X"20", X"e3", X"e3", X"20",
     X"1c", X"e2", X"08", X"8a", X"48", X"20", X"eb", X"e3",
     X"68", X"aa", X"28", X"60", X"8e", X"05", X"c0", X"48",
     X"98", X"48", X"a9", X"00", X"8d", X"fe", X"04", X"a9",
     X"07", X"8d", X"08", X"c0", X"20", X"a2", X"e2", X"f0",
     X"16", X"a8", X"6a", X"b0", X"55", X"a9", X"20", X"2c",
     X"05", X"c0", X"10", X"15", X"50", X"29", X"d0", X"4a",
     X"a9", X"10", X"2c", X"05", X"c0", X"f0", X"3b", X"a2",
     X"00", X"18", X"8e", X"fe", X"04", X"68", X"a8", X"68",
     X"60", X"98", X"29", X"18", X"f0", X"f1", X"c0", X"18",
     X"f0", X"30", X"ad", X"05", X"c0", X"c9", X"20", X"b0",
     X"29", X"c9", X"10", X"90", X"1d", X"b0", X"10", X"98",
     X"29", X"40", X"d0", X"1e", X"c0", X"10", X"90", X"12",
     X"ad", X"05", X"c0", X"29", X"10", X"d0", X"d0", X"ac",
     X"05", X"c0", X"20", X"64", X"e3", X"8c", X"05", X"c0",
     X"b0", X"05", X"ce", X"08", X"c0", X"10", X"a5", X"20",
     X"b2", X"e3", X"a2", X"01", X"38", X"b0", X"be", X"c0",
     X"20", X"b0", X"29", X"c0", X"10", X"90", X"25", X"ad",
     X"01", X"c0", X"29", X"7f", X"8d", X"13", X"03", X"4c",
     X"bc", X"e2", X"ac", X"05", X"c0", X"20", X"37", X"e3",
     X"b0", X"7b", X"a9", X"20", X"2c", X"05", X"c0", X"10",
     X"de", X"50", X"10", X"d0", X"67", X"a9", X"10", X"2c",
     X"05", X"c0", X"f0", X"2a", X"20", X"93", X"e3", X"18",
     X"58", X"90", X"fe", X"ad", X"01", X"c0", X"29", X"7f",
     X"ea", X"ea", X"cd", X"11", X"03", X"f0", X"11", X"ad",
     X"08", X"c0", X"a2", X"1c", X"20", X"1c", X"e2", X"8d",
     X"08", X"c0", X"8c", X"05", X"c0", X"b0", X"4e", X"ea",
     X"ad", X"02", X"c0", X"8d", X"12", X"03", X"98", X"29",
     X"20", X"d0", X"1a", X"20", X"93", X"e3", X"58", X"ad",
     X"18", X"03", X"30", X"fb", X"ad", X"13", X"03", X"91",
     X"fe", X"c8", X"d0", X"f3", X"e6", X"ff", X"d0", X"ef",
     X"f0", X"18", X"ea", X"ea", X"ea", X"20", X"93", X"e3",
     X"58", X"ad", X"18", X"03", X"30", X"fb", X"b1", X"fe",
     X"8d", X"13", X"03", X"c8", X"d0", X"f3", X"e6", X"ff",
     X"d0", X"ef", X"f0", X"fe", X"ad", X"05", X"c0", X"29",
     X"10", X"f0", X"c8", X"d0", X"e0", X"20", X"b2", X"e3",
     X"ad", X"fe", X"04", X"58", X"60", X"ad", X"fe", X"04",
     X"29", X"bb", X"8d", X"fe", X"04", X"58", X"60", X"ad",
     X"00", X"c0", X"29", X"03", X"aa", X"bd", X"f3", X"e3",
     X"2c", X"01", X"c0", X"10", X"02", X"09", X"10", X"8d",
     X"14", X"03", X"aa", X"ad", X"80", X"04", X"8e", X"80",
     X"04", X"29", X"7e", X"85", X"fe", X"8a", X"29", X"7e",
     X"c5", X"fe", X"f0", X"31", X"c0", X"10", X"90", X"2d",
     X"c0", X"f0", X"f0", X"29", X"ad", X"04", X"c0", X"48",
     X"a9", X"c3", X"8d", X"04", X"c0", X"ad", X"08", X"c0",
     X"a2", X"c0", X"20", X"1c", X"e2", X"8d", X"08", X"c0",
     X"68", X"8d", X"04", X"c0", X"8c", X"05", X"c0", X"ad",
     X"fe", X"04", X"d0", X"0b", X"ad", X"12", X"03", X"ea",
     X"ea", X"ea", X"8d", X"11", X"03", X"18", X"60", X"38",
     X"60", X"ea", X"ea", X"78", X"8c", X"05", X"c0", X"ad",
     X"03", X"c0", X"85", X"fe", X"ad", X"04", X"c0", X"85",
     X"ff", X"8c", X"10", X"03", X"ad", X"80", X"04", X"09",
     X"01", X"8d", X"14", X"03", X"8d", X"80", X"04", X"a0",
     X"00", X"60", X"ad", X"fe", X"04", X"a2", X"08", X"20",
     X"1c", X"e2", X"8d", X"fe", X"04", X"60", X"ea", X"ea",
     X"48", X"ad", X"14", X"03", X"30", X"19", X"68", X"ad",
     X"80", X"04", X"29", X"fe", X"8d", X"80", X"04", X"8d",
     X"14", X"03", X"68", X"68", X"68", X"ad", X"10", X"03",
     X"29", X"5d", X"8d", X"fe", X"04", X"58", X"60", X"68",
     X"4c", X"e6", X"e0", X"48", X"a9", X"40", X"8d", X"0e",
     X"03", X"68", X"60", X"48", X"a9", X"c0", X"8d", X"0e",
     X"03", X"68", X"60", X"04", X"24", X"44", X"64", X"20",
     X"06", X"e0", X"20", X"4b", X"e0", X"20", X"45", X"eb",
     X"20", X"00", X"e0", X"88", X"c8", X"20", X"60", X"e0",
     X"20", X"00", X"00", X"f0", X"55", X"c9", X"2c", X"d0",
     X"15", X"c8", X"b1", X"e9", X"c9", X"4e", X"d0", X"05",
     X"8d", X"4f", X"c1", X"10", X"e7", X"c9", X"44", X"d0",
     X"0a", X"8d", X"50", X"c1", X"10", X"de", X"a2", X"01",
     X"4c", X"1b", X"e0", X"c9", X"4a", X"d0", X"15", X"8d",
     X"41", X"c1", X"a5", X"9c", X"38", X"e9", X"02", X"8d",
     X"4d", X"c1", X"a5", X"9d", X"e9", X"00", X"8d", X"4e",
     X"c1", X"4c", X"04", X"e4", X"c9", X"41", X"d0", X"de",
     X"8d", X"4f", X"c1", X"8d", X"41", X"c1", X"c8", X"20",
     X"5d", X"e0", X"90", X"d2", X"ad", X"46", X"c1", X"8d",
     X"4e", X"c1", X"ad", X"45", X"c1", X"8d", X"4d", X"c1",
     X"b0", X"a3", X"98", X"48", X"20", X"09", X"e0", X"68",
     X"a8", X"ad", X"4c", X"c1", X"f0", X"08", X"ad", X"4f",
     X"c1", X"10", X"03", X"6c", X"4b", X"c1", X"ad", X"4b",
     X"c1", X"d0", X"03", X"4c", X"69", X"e0", X"c9", X"03",
     X"b0", X"f9", X"20", X"5a", X"e0", X"6f", X"c5", X"5f",
     X"c5", X"a5", X"92", X"85", X"9d", X"18", X"a5", X"91",
     X"69", X"02", X"85", X"9c", X"90", X"02", X"e6", X"9d",
     X"85", X"9e", X"85", X"a0", X"a5", X"9d", X"85", X"9f",
     X"85", X"a1", X"a5", X"a6", X"85", X"a2", X"a5", X"a7",
     X"85", X"a3", X"20", X"5a", X"e0", X"1f", X"c9", X"52",
     X"c9", X"20", X"5a", X"e0", X"65", X"c7", X"3a", X"c7",
     X"ad", X"4b", X"c1", X"c9", X"01", X"f0", X"08", X"2c",
     X"4f", X"c1", X"10", X"03", X"4c", X"69", X"e0", X"20",
     X"5a", X"e0", X"b5", X"c4", X"a8", X"c4", X"ad", X"2b",
     X"c1", X"8d", X"00", X"c0", X"20", X"2a", X"e0", X"20",
     X"0c", X"e0", X"e0", X"00", X"d0", X"05", X"a2", X"00",
     X"4c", X"1b", X"e0", X"bd", X"2f", X"c0", X"8d", X"01",
     X"c0", X"bd", X"2e", X"c0", X"20", X"3f", X"e8", X"a2",
     X"00", X"a0", X"02", X"10", X"02", X"8a", X"a8", X"ad",
     X"41", X"c1", X"d0", X"0c", X"b9", X"25", X"c0", X"8d",
     X"4d", X"c1", X"b9", X"26", X"c0", X"8d", X"4e", X"c1",
     X"38", X"ad", X"4d", X"c1", X"f9", X"25", X"c0", X"99",
     X"25", X"c0", X"ad", X"4e", X"c1", X"f9", X"26", X"c0",
     X"99", X"26", X"c0", X"18", X"b9", X"25", X"c0", X"79",
     X"27", X"c0", X"99", X"27", X"c0", X"b9", X"26", X"c0",
     X"79", X"28", X"c0", X"99", X"28", X"c0", X"e0", X"00",
     X"d0", X"0c", X"b9", X"2a", X"c0", X"8d", X"4c", X"c1",
     X"b9", X"29", X"c0", X"8d", X"4b", X"c1", X"ad", X"50",
     X"c1", X"30", X"36", X"ad", X"4e", X"c1", X"20", X"4d",
     X"e1", X"ad", X"4d", X"c1", X"20", X"4d", X"e1", X"a9",
     X"20", X"20", X"57", X"e0", X"b9", X"28", X"c0", X"20",
     X"4d", X"e1", X"b9", X"27", X"c0", X"20", X"4d", X"e1",
     X"ad", X"41", X"c1", X"d0", X"11", X"a9", X"20", X"20",
     X"57", X"e0", X"b9", X"2a", X"c0", X"20", X"4d", X"e1",
     X"b9", X"29", X"c0", X"20", X"4d", X"e1", X"20", X"54",
     X"e0", X"ad", X"4d", X"c1", X"85", X"0c", X"ad", X"4e",
     X"c1", X"85", X"0d", X"18", X"98", X"69", X"08", X"aa",
     X"f0", X"25", X"bd", X"23", X"c0", X"f0", X"1d", X"c9",
     X"ff", X"d0", X"03", X"4c", X"f5", X"e4", X"8d", X"41",
     X"c1", X"a0", X"00", X"e8", X"bd", X"23", X"c0", X"91",
     X"0c", X"e6", X"0c", X"d0", X"02", X"e6", X"0d", X"ce",
     X"41", X"c1", X"d0", X"ef", X"e8", X"d0", X"db", X"ad",
     X"23", X"c0", X"8d", X"01", X"c0", X"ad", X"24", X"c0",
     X"f0", X"07", X"20", X"3f", X"e8", X"a2", X"02", X"10",
     X"c9", X"60", X"a9", X"ff", X"8d", X"4f", X"c1", X"8d",
     X"50", X"c1", X"8d", X"3c", X"c1", X"a9", X"00", X"8d",
     X"4d", X"c1", X"8d", X"4e", X"c1", X"8d", X"41", X"c1",
     X"60", X"46", X"69", X"6c", X"65", X"20", X"6e", X"6f",
     X"74", X"20", X"66", X"6f", X"75", X"6e", X"64", X"00",
     X"49", X"6e", X"76", X"61", X"6c", X"69", X"64", X"20",
     X"63", X"6f", X"6d", X"6d", X"61", X"6e", X"64", X"20",
     X"65", X"6e", X"64", X"00", X"4e", X"6f", X"20", X"64",
     X"72", X"69", X"76", X"65", X"20", X"6e", X"75", X"6d",
     X"62", X"65", X"72", X"00", X"42", X"61", X"64", X"20",
     X"64", X"72", X"69", X"76", X"65", X"20", X"6e", X"75",
     X"6d", X"62", X"65", X"72", X"00", X"49", X"6e", X"76",
     X"61", X"6c", X"69", X"64", X"20", X"66", X"69", X"6c",
     X"65", X"6e", X"61", X"6d", X"65", X"00", X"44", X"69",
     X"73", X"63", X"20", X"65", X"72", X"72", X"6f", X"72",
     X"00", X"49", X"6c", X"6c", X"65", X"67", X"61", X"6c",
     X"20", X"61", X"74", X"74", X"72", X"69", X"62", X"75",
     X"74", X"65", X"00", X"57", X"69", X"6c", X"64", X"63",
     X"61", X"72", X"64", X"28", X"73", X"29", X"20", X"6e",
     X"6f", X"74", X"20", X"61", X"6c", X"6c", X"6f", X"77",
     X"65", X"64", X"00", X"46", X"69", X"6c", X"65", X"20",
     X"61", X"6c", X"72", X"65", X"61", X"64", X"79", X"20",
     X"65", X"78", X"69", X"73", X"74", X"73", X"00", X"49",
     X"6e", X"73", X"75", X"66", X"66", X"69", X"63", X"69",
     X"65", X"6e", X"74", X"20", X"64", X"69", X"73", X"6b",
     X"20", X"73", X"70", X"61", X"63", X"65", X"00", X"53",
     X"74", X"61", X"72", X"74", X"20", X"61", X"64", X"64",
     X"72", X"65", X"73", X"73", X"20", X"6d", X"69", X"73",
     X"73", X"69", X"6e", X"67", X"00", X"49", X"6c", X"6c",
     X"65", X"67", X"61", X"6c", X"20", X"71", X"75", X"61",
     X"6e", X"74", X"69", X"74", X"79", X"00", X"45", X"6e",
     X"64", X"20", X"61", X"64", X"64", X"72", X"65", X"73",
     X"73", X"20", X"6d", X"69", X"73", X"73", X"69", X"6e",
     X"67", X"00", X"53", X"74", X"61", X"72", X"74", X"20",
     X"61", X"64", X"64", X"72", X"65", X"73", X"73", X"20",
     X"3e", X"20", X"65", X"6e", X"64", X"20", X"61", X"64",
     X"64", X"72", X"65", X"73", X"73", X"00", X"4d", X"69",
     X"73", X"73", X"69", X"6e", X"67", X"20", X"27", X"54",
     X"4f", X"27", X"00", X"52", X"65", X"6e", X"61", X"6d",
     X"65", X"64", X"20", X"66", X"69", X"6c", X"65", X"20",
     X"6e", X"6f", X"74", X"20", X"6f", X"6e", X"20", X"73",
     X"61", X"6d", X"65", X"20", X"64", X"69", X"73", X"6b",
     X"00", X"4d", X"69", X"73", X"73", X"69", X"6e", X"67",
     X"20", X"63", X"6f", X"6d", X"6d", X"61", X"00", X"53",
     X"6f", X"75", X"72", X"63", X"65", X"20", X"61", X"6e",
     X"64", X"20", X"64", X"65", X"73", X"74", X"69", X"6e",
     X"61", X"74", X"69", X"6f", X"6e", X"20", X"64", X"72",
     X"69", X"76", X"65", X"73", X"20", X"6d", X"75", X"73",
     X"74", X"20", X"62", X"65", X"20", X"73", X"61", X"6d",
     X"65", X"00", X"44", X"65", X"73", X"74", X"69", X"6e",
     X"61", X"74", X"69", X"6f", X"6e", X"20", X"6e", X"6f",
     X"74", X"20", X"73", X"70", X"65", X"63", X"69", X"66",
     X"69", X"65", X"64", X"00", X"43", X"61", X"6e", X"6e",
     X"6f", X"74", X"20", X"6d", X"65", X"72", X"67", X"65",
     X"20", X"61", X"6e", X"64", X"20", X"6f", X"76", X"65",
     X"72", X"77", X"72", X"69", X"74", X"65", X"00", X"53",
     X"69", X"6e", X"67", X"6c", X"65", X"20", X"64", X"65",
     X"73", X"74", X"69", X"6e", X"61", X"74", X"69", X"6f",
     X"6e", X"20", X"66", X"69", X"6c", X"65", X"20", X"6e",
     X"6f", X"74", X"20", X"61", X"6c", X"6c", X"6f", X"77",
     X"65", X"64", X"00", X"53", X"79", X"6e", X"74", X"61",
     X"78", X"20", X"65", X"72", X"72", X"6f", X"72", X"00",
     X"d9", X"e8", X"fc", X"0c", X"1d", X"2e", X"39", X"4b",
     X"63", X"77", X"8f", X"a5", X"b6", X"ca", X"e6", X"f3",
     X"11", X"1f", X"4a", X"64", X"7f", X"a3", X"e5", X"e5",
     X"e5", X"e6", X"e6", X"e6", X"e6", X"e6", X"e6", X"e6",
     X"e6", X"e6", X"e6", X"e6", X"e6", X"e6", X"e7", X"e7",
     X"e7", X"e7", X"e7", X"e7", X"e8", X"8e", X"ff", X"04",
     X"6c", X"49", X"c1", X"ca", X"ad", X"fd", X"04", X"29",
     X"01", X"f0", X"03", X"4c", X"69", X"e0", X"e0", X"16",
     X"b0", X"15", X"bd", X"b0", X"e7", X"85", X"0c", X"bd",
     X"c6", X"e7", X"85", X"0d", X"20", X"2d", X"e0", X"a9",
     X"3a", X"20", X"57", X"e0", X"4c", X"13", X"e8", X"8a",
     X"20", X"4d", X"e1", X"ad", X"fe", X"04", X"f0", X"03",
     X"20", X"4d", X"e1", X"4c", X"ff", X"e1", X"60", X"20",
     X"06", X"e2", X"ad", X"fe", X"04", X"f0", X"05", X"a2",
     X"05", X"4c", X"1b", X"e0", X"60", X"20", X"0a", X"e2",
     X"4c", X"1a", X"e8", X"a9", X"23", X"8d", X"03", X"c0",
     X"a9", X"c0", X"8d", X"04", X"c0", X"a9", X"00", X"8d",
     X"01", X"c0", X"8d", X"0a", X"c0", X"a9", X"01", X"8d",
     X"02", X"c0", X"20", X"24", X"e0", X"60", X"ae", X"00",
     X"c0", X"bd", X"13", X"c0", X"f0", X"01", X"60", X"a2",
     X"03", X"4c", X"1b", X"e0", X"a0", X"00", X"b1", X"0c",
     X"f0", X"06", X"20", X"57", X"e0", X"c8", X"10", X"f6",
     X"60", X"ad", X"46", X"c1", X"d0", X"09", X"ad", X"45",
     X"c1", X"30", X"04", X"c9", X"04", X"30", X"02", X"a9",
     X"ff", X"60", X"20", X"27", X"e0", X"a2", X"07", X"bd",
     X"33", X"c0", X"9d", X"23", X"c1", X"ca", X"10", X"f7",
     X"60", X"20", X"27", X"e0", X"a2", X"07", X"bd", X"23",
     X"c1", X"9d", X"33", X"c0", X"ca", X"10", X"f7", X"20",
     X"21", X"e0", X"60", X"ad", X"3e", X"c1", X"8d", X"01",
     X"c0", X"ad", X"3d", X"c1", X"20", X"3f", X"e8", X"a2",
     X"00", X"ac", X"3f", X"c1", X"bd", X"2c", X"c1", X"99",
     X"23", X"c0", X"c8", X"e8", X"e0", X"10", X"d0", X"f4",
     X"ee", X"25", X"c0", X"20", X"21", X"e0", X"60", X"20",
     X"3f", X"e0", X"f0", X"08", X"ee", X"29", X"c1", X"d0",
     X"03", X"ee", X"2a", X"c1", X"60", X"ad", X"23", X"c1",
     X"f0", X"2b", X"8d", X"02", X"c0", X"ad", X"24", X"c1",
     X"8d", X"01", X"c0", X"20", X"24", X"e0", X"ad", X"24",
     X"c0", X"8d", X"23", X"c1", X"ad", X"23", X"c0", X"8d",
     X"24", X"c1", X"38", X"ad", X"27", X"c1", X"e9", X"01",
     X"8d", X"27", X"c1", X"ad", X"28", X"c1", X"e9", X"00",
     X"8d", X"28", X"c1", X"a9", X"01", X"60", X"20", X"24",
     X"e0", X"ad", X"25", X"c0", X"c9", X"0f", X"d0", X"31",
     X"ad", X"24", X"c0", X"f0", X"0c", X"8d", X"02", X"c0",
     X"ad", X"23", X"c0", X"8d", X"01", X"c0", X"4c", X"f6",
     X"e8", X"ad", X"23", X"c1", X"f0", X"39", X"8d", X"24",
     X"c0", X"ad", X"24", X"c1", X"8d", X"23", X"c0", X"20",
     X"21", X"e0", X"20", X"3f", X"e0", X"a9", X"00", X"aa",
     X"9d", X"23", X"c0", X"e8", X"d0", X"fa", X"20", X"21",
     X"e0", X"a2", X"03", X"bd", X"23", X"c0", X"f0", X"07",
     X"8a", X"18", X"69", X"10", X"aa", X"d0", X"f4", X"8a",
     X"8d", X"3f", X"c1", X"ad", X"01", X"c0", X"8d", X"3e",
     X"c1", X"ad", X"02", X"c0", X"8d", X"3d", X"c1", X"60",
     X"20", X"24", X"e0", X"ae", X"3f", X"c1", X"d0", X"28",
     X"20", X"24", X"e0", X"a2", X"03", X"a9", X"26", X"85",
     X"0c", X"a9", X"c0", X"85", X"0d", X"a0", X"00", X"b1",
     X"0c", X"f0", X"15", X"a0", X"08", X"b9", X"2c", X"c1",
     X"c9", X"3f", X"f0", X"04", X"d1", X"0c", X"d0", X"08",
     X"88", X"10", X"f2", X"8a", X"8d", X"3f", X"c1", X"60",
     X"8a", X"18", X"69", X"10", X"b0", X"0e", X"aa", X"a5",
     X"0c", X"69", X"10", X"85", X"0c", X"90", X"d6", X"e6",
     X"0d", X"4c", X"65", X"e9", X"ad", X"24", X"c0", X"f0",
     X"0c", X"8d", X"02", X"c0", X"ad", X"23", X"c0", X"8d",
     X"01", X"c0", X"4c", X"58", X"e9", X"a2", X"00", X"60",
     X"ad", X"13", X"c0", X"d0", X"fa", X"8d", X"00", X"c0",
     X"a9", X"13", X"8d", X"03", X"c0", X"a9", X"c0", X"8d",
     X"04", X"c0", X"4c", X"35", X"e8", X"20", X"20", X"20",
     X"20", X"20", X"20", X"20", X"20", X"20", X"20", X"20",
     X"20", X"00", X"a2", X"0b", X"a9", X"20", X"9d", X"bd",
     X"e9", X"ca", X"10", X"fa", X"20", X"60", X"e0", X"20",
     X"00", X"00", X"f0", X"69", X"38", X"e9", X"30", X"c9",
     X"04", X"b0", X"0f", X"c8", X"8d", X"2b", X"c1", X"a2",
     X"09", X"a9", X"20", X"9d", X"2b", X"c1", X"ca", X"d0",
     X"fa", X"60", X"a5", X"ea", X"48", X"a5", X"e9", X"48",
     X"98", X"18", X"65", X"e9", X"85", X"e9", X"90", X"02",
     X"e6", X"ea", X"20", X"5a", X"e0", X"8b", X"ce", X"17",
     X"cf", X"24", X"28", X"10", X"56", X"20", X"5a", X"e0",
     X"15", X"d7", X"d0", X"d7", X"c9", X"0c", X"90", X"02",
     X"a9", X"0c", X"a8", X"88", X"30", X"08", X"b1", X"91",
     X"99", X"bd", X"e9", X"4c", X"1b", X"ea", X"a5", X"e9",
     X"48", X"a9", X"bd", X"85", X"e9", X"a9", X"e9", X"85",
     X"ea", X"c8", X"20", X"45", X"ea", X"68", X"85", X"ea",
     X"68", X"18", X"85", X"e9", X"e5", X"ea", X"49", X"ff",
     X"a8", X"68", X"85", X"ea", X"60", X"ad", X"0c", X"c0",
     X"8d", X"2b", X"c1", X"20", X"e7", X"e9", X"c8", X"b1",
     X"e9", X"88", X"c9", X"cd", X"f0", X"04", X"c9", X"2d",
     X"d0", X"13", X"b1", X"e9", X"38", X"e9", X"30", X"c9",
     X"04", X"90", X"05", X"a2", X"04", X"4c", X"1b", X"e0",
     X"8d", X"2b", X"c1", X"c8", X"c8", X"a2", X"00", X"a9",
     X"06", X"20", X"8c", X"ea", X"b1", X"e9", X"c9", X"2e",
     X"d0", X"08", X"c8", X"a2", X"06", X"a9", X"03", X"20",
     X"8c", X"ea", X"20", X"00", X"00", X"f0", X"04", X"c9",
     X"20", X"d0", X"d8", X"60", X"8d", X"41", X"c1", X"b1",
     X"e9", X"c9", X"2a", X"f0", X"16", X"c9", X"3f", X"f0",
     X"07", X"20", X"4e", X"e0", X"c9", X"00", X"f0", X"0a",
     X"9d", X"2c", X"c1", X"e8", X"c8", X"ce", X"41", X"c1",
     X"d0", X"e5", X"60", X"a9", X"3f", X"9d", X"2c", X"c1",
     X"e8", X"ce", X"41", X"c1", X"d0", X"f7", X"c8", X"60",
     X"c9", X"30", X"90", X"14", X"c9", X"3a", X"90", X"12",
     X"c9", X"41", X"90", X"0c", X"c9", X"5b", X"90", X"0a",
     X"c9", X"61", X"90", X"04", X"c9", X"7b", X"90", X"02",
     X"a9", X"00", X"60", X"20", X"33", X"e0", X"ad", X"26",
     X"c1", X"8d", X"01", X"c0", X"ad", X"25", X"c1", X"8d",
     X"02", X"c0", X"a9", X"00", X"8d", X"3f", X"c1", X"4c",
     X"45", X"e0", X"a2", X"09", X"ac", X"3f", X"c1", X"b9",
     X"2c", X"c0", X"9d", X"2c", X"c1", X"c8", X"e8", X"e0",
     X"10", X"d0", X"f4", X"60", X"ae", X"3f", X"c1", X"a0",
     X"06", X"bd", X"23", X"c0", X"c9", X"20", X"d0", X"03",
     X"20", X"57", X"e0", X"e8", X"88", X"d0", X"f2", X"ae",
     X"3f", X"c1", X"a0", X"06", X"bd", X"23", X"c0", X"c9",
     X"20", X"f0", X"03", X"20", X"57", X"e0", X"e8", X"88",
     X"d0", X"f2", X"a9", X"2e", X"20", X"57", X"e0", X"a0",
     X"03", X"bd", X"23", X"c0", X"20", X"57", X"e0", X"e8",
     X"88", X"d0", X"f6", X"60", X"a5", X"0c", X"8d", X"47",
     X"c1", X"a5", X"0d", X"8d", X"48", X"c1", X"ba", X"e8",
     X"e8", X"8e", X"40", X"c1", X"60", X"a2", X"08", X"bd",
     X"2c", X"c1", X"c9", X"3f", X"f0", X"2b", X"ca", X"10",
     X"f6", X"60", X"43", X"4f", X"4d", X"20", X"06", X"e0",
     X"a0", X"00", X"98", X"20", X"48", X"ea", X"ad", X"32",
     X"c1", X"c9", X"20", X"d0", X"0b", X"a2", X"02", X"bd",
     X"52", X"eb", X"9d", X"32", X"c1", X"ca", X"10", X"f7",
     X"20", X"45", X"eb", X"20", X"00", X"e0", X"4c", X"62",
     X"e4", X"a2", X"07", X"4c", X"1b", X"e0", X"78", X"d8",
     X"a2", X"ff", X"9a", X"e8", X"8a", X"a8", X"ca", X"d0",
     X"fd", X"88", X"d0", X"fa", X"9d", X"00", X"c0", X"9d",
     X"00", X"c1", X"95", X"00", X"9d", X"00", X"02", X"ca",
     X"d0", X"f2", X"a2", X"7a", X"bd", X"ed", X"ee", X"9d",
     X"80", X"04", X"ca", X"10", X"f7", X"20", X"ae", X"ee",
     X"a2", X"0c", X"bd", X"68", X"ef", X"9d", X"e0", X"bf",
     X"ca", X"10", X"f7", X"20", X"e0", X"bf", X"c0", X"ea",
     X"f0", X"0f", X"a9", X"01", X"8d", X"07", X"c0", X"a9",
     X"44", X"8d", X"dc", X"04", X"a9", X"47", X"8d", X"e4",
     X"04", X"a2", X"ff", X"86", X"a9", X"a9", X"ff", X"a0",
     X"97", X"85", X"a6", X"84", X"a7", X"8d", X"c1", X"02",
     X"8c", X"c2", X"02", X"85", X"a2", X"84", X"a3", X"a2",
     X"1c", X"bd", X"cf", X"ee", X"95", X"e1", X"ca", X"d0",
     X"f8", X"ad", X"07", X"c0", X"f0", X"28", X"a9", X"b9",
     X"85", X"f0", X"a9", X"ec", X"85", X"f1", X"a9", X"20",
     X"8d", X"4e", X"02", X"a9", X"04", X"8d", X"4f", X"02",
     X"a9", X"00", X"8d", X"60", X"02", X"a2", X"12", X"bd",
     X"5d", X"ee", X"9d", X"38", X"02", X"ca", X"10", X"f7",
     X"a9", X"b0", X"a0", X"cc", X"30", X"19", X"a9", X"ff",
     X"a0", X"bf", X"8d", X"e1", X"02", X"8c", X"e2", X"02",
     X"a2", X"08", X"bd", X"54", X"ee", X"9d", X"28", X"02",
     X"ca", X"10", X"f7", X"a9", X"ed", X"a0", X"cb", X"85",
     X"1b", X"84", X"1c", X"a9", X"4c", X"85", X"1a", X"85",
     X"c3", X"85", X"21", X"8d", X"fb", X"02", X"a9", X"a0",
     X"a0", X"d2", X"ae", X"07", X"c0", X"f0", X"04", X"a9",
     X"36", X"a0", X"d3", X"85", X"22", X"84", X"23", X"8d",
     X"fc", X"02", X"8c", X"fd", X"02", X"a9", X"c4", X"a0",
     X"04", X"8d", X"f5", X"02", X"8c", X"f6", X"02", X"a9",
     X"00", X"8d", X"ff", X"04", X"8d", X"fd", X"04", X"20",
     X"5a", X"e0", X"88", X"f8", X"b8", X"f8", X"a9", X"50",
     X"85", X"31", X"a9", X"30", X"85", X"32", X"a9", X"03",
     X"85", X"c2", X"a9", X"00", X"85", X"d7", X"85", X"88",
     X"85", X"2f", X"48", X"8d", X"00", X"05", X"8d", X"01",
     X"05", X"8d", X"02", X"05", X"8d", X"f7", X"02", X"85",
     X"2e", X"8d", X"f1", X"02", X"8d", X"f2", X"02", X"8d",
     X"f4", X"02", X"a9", X"88", X"85", X"85", X"a9", X"02",
     X"8d", X"c0", X"02", X"a9", X"01", X"a0", X"05", X"85",
     X"9a", X"84", X"9b", X"a9", X"03", X"85", X"9c", X"84",
     X"9d", X"85", X"9e", X"84", X"9f", X"85", X"a0", X"84",
     X"a1", X"a2", X"00", X"20", X"92", X"ee", X"a2", X"09",
     X"bd", X"40", X"ee", X"9d", X"2b", X"c1", X"ca", X"10",
     X"f7", X"a9", X"8a", X"8d", X"49", X"c1", X"a9", X"ee",
     X"8d", X"4a", X"c1", X"a2", X"d8", X"8e", X"10", X"03",
     X"a2", X"08", X"20", X"03", X"e0", X"20", X"48", X"e0",
     X"20", X"00", X"e0", X"20", X"09", X"e0", X"20", X"a3",
     X"ee", X"a2", X"08", X"bd", X"5a", X"ed", X"95", X"35",
     X"ca", X"10", X"f8", X"a2", X"ff", X"e8", X"bd", X"d0",
     X"9f", X"9d", X"82", X"bb", X"d0", X"f7", X"a2", X"1a",
     X"bd", X"3f", X"ed", X"9d", X"e0", X"bf", X"ca", X"10",
     X"f7", X"a9", X"ae", X"a0", X"ed", X"ae", X"07", X"c0",
     X"f0", X"04", X"a9", X"f1", X"a0", X"ed", X"85", X"0c",
     X"84", X"0d", X"20", X"2d", X"e0", X"a2", X"09", X"bd",
     X"4a", X"ee", X"9d", X"2b", X"c1", X"ca", X"10", X"f7",
     X"20", X"0c", X"e0", X"e0", X"00", X"d0", X"0d", X"86",
     X"35", X"a9", X"35", X"85", X"0c", X"a9", X"ee", X"85",
     X"0d", X"20", X"2d", X"e0", X"4c", X"e0", X"bf", X"78",
     X"a9", X"84", X"8d", X"80", X"04", X"8d", X"14", X"03",
     X"20", X"f8", X"bf", X"a2", X"34", X"a0", X"00", X"58",
     X"20", X"5a", X"d4", X"cd", X"c4", X"bd", X"c4", X"6c",
     X"4b", X"c1", X"21", X"42", X"4f", X"4f", X"54", X"55",
     X"50", X"00", X"00", X"69", X"6e", X"73", X"65", X"72",
     X"74", X"20", X"73", X"79", X"73", X"74", X"65", X"6d",
     X"20", X"64", X"69", X"73", X"63", X"00", X"0c", X"4e",
     X"6f", X"20", X"6f", X"70", X"65", X"72", X"61", X"74",
     X"69", X"6e", X"67", X"20", X"73", X"79", X"73", X"74",
     X"65", X"6d", X"20", X"6f", X"6e", X"20", X"64", X"69",
     X"73", X"63", X"08", X"00", X"0c", X"52", X"56", X"31",
     X"20", X"61", X"64", X"6a", X"75", X"73", X"74", X"6d",
     X"65", X"6e", X"74", X"20", X"72", X"65", X"71", X"75",
     X"69", X"72", X"65", X"64", X"08", X"00", X"0c", X"4f",
     X"52", X"49", X"43", X"20", X"45", X"58", X"54", X"45",
     X"4e", X"44", X"45", X"44", X"20", X"42", X"41", X"53",
     X"49", X"43", X"20", X"56", X"31", X"2e", X"30", X"0d",
     X"0a", X"60", X"20", X"31", X"39", X"38", X"33", X"20",
     X"54", X"41", X"4e", X"47", X"45", X"52", X"49", X"4e",
     X"45", X"0d", X"0a", X"0a", X"0a", X"34", X"37", X"38",
     X"37", X"30", X"20", X"42", X"59", X"54", X"45", X"53",
     X"20", X"46", X"52", X"45", X"45", X"0d", X"0a", X"0a",
     X"00", X"0c", X"4f", X"52", X"49", X"43", X"20", X"45",
     X"58", X"54", X"45", X"4e", X"44", X"45", X"44", X"20",
     X"42", X"41", X"53", X"49", X"43", X"20", X"56", X"31",
     X"2e", X"31", X"0d", X"0a", X"60", X"20", X"31", X"39",
     X"38", X"33", X"20", X"54", X"41", X"4e", X"47", X"45",
     X"52", X"49", X"4e", X"45", X"0d", X"0a", X"0a", X"0a",
     X"20", X"33", X"37", X"36", X"33", X"31", X"20", X"42",
     X"59", X"54", X"45", X"53", X"20", X"46", X"52", X"45",
     X"45", X"0d", X"0a", X"0a", X"00", X"0d", X"0a", X"52",
     X"65", X"61", X"64", X"79", X"20", X"0d", X"0a", X"00",
     X"00", X"53", X"59", X"53", X"54", X"45", X"4d", X"44",
     X"4f", X"53", X"00", X"42", X"4f", X"4f", X"54", X"55",
     X"50", X"43", X"4f", X"4d", X"4c", X"03", X"ec", X"4c",
     X"30", X"f4", X"01", X"00", X"40", X"4c", X"7c", X"f7",
     X"4c", X"78", X"eb", X"4c", X"c1", X"f5", X"4c", X"65",
     X"f8", X"4c", X"22", X"ee", X"4c", X"b2", X"f8", X"40",
     X"a2", X"31", X"a0", X"00", X"a9", X"1a", X"99", X"80",
     X"bb", X"99", X"80", X"bc", X"99", X"80", X"bd", X"99",
     X"80", X"be", X"99", X"fe", X"be", X"88", X"d0", X"ee",
     X"f0", X"02", X"a2", X"13", X"20", X"92", X"ee", X"4c",
     X"8f", X"ee", X"20", X"a3", X"ee", X"4c", X"9d", X"ee",
     X"e8", X"99", X"82", X"bb", X"c8", X"bd", X"63", X"ed",
     X"d0", X"f6", X"60", X"a0", X"1b", X"a9", X"20", X"99",
     X"81", X"bb", X"88", X"d0", X"fa", X"60", X"a2", X"00",
     X"bd", X"a5", X"c0", X"a8", X"a9", X"55", X"9d", X"a5",
     X"c0", X"dd", X"a5", X"c0", X"d0", X"b2", X"a9", X"aa",
     X"9d", X"a5", X"c0", X"dd", X"a5", X"c0", X"d0", X"a8",
     X"98", X"9d", X"a5", X"c0", X"e8", X"d0", X"e1", X"60",
     X"e6", X"e9", X"d0", X"02", X"e6", X"ea", X"ad", X"60",
     X"ea", X"c9", X"20", X"f0", X"f3", X"20", X"41", X"ea",
     X"60", X"2c", X"60", X"ea", X"2c", X"60", X"ea", X"60",
     X"80", X"4f", X"c7", X"52", X"58", X"04", X"00", X"00",
     X"00", X"4c", X"60", X"ea", X"4c", X"e6", X"04", X"4c",
     X"d6", X"04", X"4c", X"de", X"04", X"08", X"78", X"8d",
     X"82", X"04", X"68", X"8d", X"83", X"04", X"ad", X"80",
     X"04", X"48", X"ad", X"81", X"04", X"20", X"e6", X"04",
     X"ad", X"83", X"04", X"48", X"ad", X"82", X"04", X"28",
     X"20", X"84", X"04", X"08", X"78", X"8d", X"82", X"04",
     X"68", X"8d", X"83", X"04", X"68", X"20", X"e6", X"04",
     X"ad", X"83", X"04", X"48", X"ad", X"82", X"04", X"28",
     X"60", X"a9", X"00", X"8d", X"81", X"04", X"a9", X"66",
     X"8d", X"85", X"04", X"a9", X"d4", X"8d", X"86", X"04",
     X"4c", X"90", X"04", X"08", X"ba", X"fe", X"02", X"01",
     X"4c", X"28", X"02", X"08", X"ba", X"fe", X"02", X"01",
     X"4c", X"2b", X"02", X"78", X"29", X"02", X"8d", X"81",
     X"04", X"ad", X"80", X"04", X"29", X"fd", X"0d", X"81",
     X"04", X"8d", X"14", X"03", X"8d", X"80", X"04", X"60",
     X"a9", X"06", X"20", X"87", X"04", X"ac", X"02", X"c0",
     X"a9", X"00", X"4c", X"87", X"04", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff", X"ff",
     X"4f", X"72", X"69", X"63", X"20", X"44", X"4f", X"53",
     X"20", X"56", X"30", X"2e", X"36", X"00", X"00", X"00",
     X"28", X"43", X"29", X"20", X"4f", X"52", X"49", X"43",
     X"20", X"31", X"39", X"38", X"33", X"00", X"00", X"00",
     X"00", X"00", X"00", X"00", X"00", X"00", X"00", X"00",
     X"00", X"00", X"ae", X"e0", X"7e", X"eb", X"c0", X"e3");

begin

process (clk)
  begin
    if rising_edge(clk) then
      data <= rom_data(TO_INTEGER(unsigned(addr)));
    end if;
  end process;

end architecture;
